
module BP_NB32_BP_LEN4_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   net409532, net409531, net409506, net409505, net409501, net409498,
         net409494, net409493, net409490, net409484, net409481, net409480,
         net409479, net409478, net409475, net409474, net409473, net409471,
         net409470, net409469, net409468, net409467, net409466, net409465,
         net409463, net409461, net409460, net409457, net409455, net409442,
         net409438, net409431, net409426, net409425, net409424, net409423,
         net409422, net409421, net409420, net409419, net409416, net409412,
         net409410, net409407, net409403, net409402, net409401, net409400,
         net409399, net409398, net409397, net409383, net409382, net409380,
         net409375, net409368, net409363, net409358, net409357, net409352,
         net409351, net409346, net409338, net409325, net409324, net409323,
         net409322, net409320, net409318, net409317, net409316, net409315,
         net409313, net409312, net409310, net409309, net409308, net409305,
         net409304, net409302, net409301, net409300, net409299, net409298,
         net409295, net409294, net412778, net412777, net412793, net412803,
         net412807, net412813, net412837, net412839, net412841, net412844,
         net412845, net412849, net412854, net412864, net412863, net409328,
         net409327, net421184, net412835, net412826, net421857, net421917,
         net421916, net421914, net422133, net422142, net422148, net422152,
         net422154, net422162, net422175, net409321, net424932, net424910,
         net409365, net409364, net409362, net425779, net425902, net425903,
         net425890, net425889, net425863, net425858, net425847, net409319,
         net409311, net409303, net421930, net421921, net422158, net409451,
         net409450, net412860, net409495, net409488, net409487, net409486,
         net409464, net409462, net409459, net409458, net409456, net409454,
         net409453, net409452, net409449, net409448, net409447, net409446,
         net425920, net424880, net409394, net409393, net409392, net409391,
         net409390, net409355, net409353, net424929, net424928, net424911,
         net424901, net424887, net424869, net424868, net424857, net422128,
         net412829, net409418, net409395, net425918, net412858, net412825,
         net412819, net409520, net409514, net409513, net409512, net409511,
         net409307, net409306, net409297, net421923, net421879, net409359,
         net409354, net409350, net409349, net409348, net421936, net421933,
         net421877, net409356, net409337, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85;

  NAND4_X2 net425791 ( .A1(net425863), .A2(net425858), .A3(net409362), .A4(
        net409363), .ZN(net409351) );
  NAND2_X2 net409374 ( .A1(net409362), .A2(n29), .ZN(net422133) );
  NAND2_X2 net425807 ( .A1(net409362), .A2(net409365), .ZN(net409380) );
  NAND2_X2 net425809 ( .A1(net409363), .A2(net409364), .ZN(net409383) );
  NAND2_X2 net425808 ( .A1(net421857), .A2(net409364), .ZN(net409382) );
  NAND2_X2 net425795 ( .A1(n17), .A2(net409364), .ZN(net409355) );
  NAND3_X1 syn233 ( .A1(net412849), .A2(net409391), .A3(net409392), .ZN(
        net424869) );
  AND2_X2 syn115 ( .A1(net409393), .A2(net409391), .ZN(n11) );
  INV_X2 net425832 ( .A(B[31]), .ZN(net422175) );
  INV_X2 net421855 ( .A(A[29]), .ZN(net409356) );
  NAND2_X1 U2 ( .A1(net421933), .A2(n2), .ZN(n3) );
  XNOR2_X1 U3 ( .A(n3), .B(net421930), .ZN(SUM[30]) );
  NAND2_X1 U4 ( .A1(net421936), .A2(net409337), .ZN(net421933) );
  NAND2_X1 U5 ( .A1(net425779), .A2(A[29]), .ZN(n2) );
  AND2_X1 U6 ( .A1(net421921), .A2(n2), .ZN(net421916) );
  BUF_X4 U7 ( .A(B[31]), .Z(net425779) );
  NAND2_X1 U8 ( .A1(net421879), .A2(net409349), .ZN(net421936) );
  CLKBUF_X1 U9 ( .A(net421936), .Z(net412793) );
  NAND2_X1 U10 ( .A1(net422175), .A2(net409356), .ZN(net409337) );
  NAND2_X1 U11 ( .A1(net409337), .A2(n1), .ZN(net409346) );
  NAND2_X1 U12 ( .A1(net421877), .A2(net409337), .ZN(net421917) );
  NAND2_X1 U13 ( .A1(net425779), .A2(A[29]), .ZN(n1) );
  NAND2_X1 U14 ( .A1(net421879), .A2(net409349), .ZN(net421877) );
  NAND2_X1 U15 ( .A1(net424887), .A2(net421923), .ZN(net421879) );
  INV_X1 U16 ( .A(net409348), .ZN(net421923) );
  NAND2_X1 U17 ( .A1(net409353), .A2(net409354), .ZN(net409348) );
  INV_X1 U18 ( .A(net409355), .ZN(net409354) );
  NOR2_X2 U19 ( .A1(net409350), .A2(net409351), .ZN(net409349) );
  INV_X1 U20 ( .A(net409352), .ZN(net409350) );
  BUF_X1 U21 ( .A(net424887), .Z(net421857) );
  NAND2_X1 U22 ( .A1(net409352), .A2(net409353), .ZN(net409357) );
  OAI21_X1 U23 ( .B1(net412835), .B2(net409355), .A(net409359), .ZN(net409358)
         );
  INV_X1 U24 ( .A(net409351), .ZN(net409359) );
  NAND2_X1 U25 ( .A1(net412825), .A2(net409511), .ZN(net409297) );
  CLKBUF_X1 U26 ( .A(net409297), .Z(net412841) );
  NAND3_X1 U27 ( .A1(net409297), .A2(net409449), .A3(net409448), .ZN(net409447) );
  NOR2_X1 U28 ( .A1(net409514), .A2(net409513), .ZN(net412825) );
  NAND3_X1 U29 ( .A1(net409324), .A2(net412819), .A3(net409323), .ZN(net409511) );
  AND2_X1 U30 ( .A1(net409512), .A2(net409511), .ZN(net412803) );
  AND4_X1 U31 ( .A1(net409318), .A2(net412858), .A3(net409304), .A4(net425918), 
        .ZN(net412819) );
  CLKBUF_X1 U32 ( .A(net409319), .Z(net412858) );
  INV_X1 U33 ( .A(net412858), .ZN(net409310) );
  OAI21_X1 U34 ( .B1(n4), .B2(n5), .A(net409307), .ZN(net409514) );
  NOR2_X1 U35 ( .A1(net409513), .A2(net409514), .ZN(net409512) );
  NAND2_X1 U36 ( .A1(net409304), .A2(n10), .ZN(n5) );
  OR2_X1 U37 ( .A1(B[7]), .A2(A[7]), .ZN(n10) );
  AND2_X1 U38 ( .A1(n7), .A2(n8), .ZN(n4) );
  AND2_X1 U39 ( .A1(net409303), .A2(net409311), .ZN(n8) );
  NAND2_X1 U40 ( .A1(net409319), .A2(n6), .ZN(n7) );
  AND2_X1 U41 ( .A1(B[4]), .A2(A[4]), .ZN(n6) );
  NOR2_X1 U42 ( .A1(net409520), .A2(net409322), .ZN(net409513) );
  NAND4_X1 U43 ( .A1(net409318), .A2(net409319), .A3(net409304), .A4(net409306), .ZN(net409520) );
  OR2_X1 U44 ( .A1(B[7]), .A2(A[7]), .ZN(net409306) );
  NAND2_X1 U45 ( .A1(net409323), .A2(net409324), .ZN(net409321) );
  NAND2_X2 U46 ( .A1(net409322), .A2(net409324), .ZN(net409325) );
  CLKBUF_X1 U47 ( .A(net409323), .Z(net412864) );
  NAND2_X1 U48 ( .A1(net425918), .A2(net409307), .ZN(net409300) );
  CLKBUF_X1 U49 ( .A(B[7]), .Z(n9) );
  OR2_X1 U50 ( .A1(B[7]), .A2(A[7]), .ZN(net425918) );
  NAND2_X1 U51 ( .A1(n9), .A2(A[7]), .ZN(net409307) );
  NAND2_X1 U52 ( .A1(net409302), .A2(net409303), .ZN(net409301) );
  NAND2_X1 U53 ( .A1(net409304), .A2(net409303), .ZN(net409308) );
  OAI21_X2 U54 ( .B1(net409309), .B2(net409310), .A(net409311), .ZN(net409305)
         );
  NAND2_X1 U55 ( .A1(net422128), .A2(net424928), .ZN(net424887) );
  NAND2_X1 U56 ( .A1(net424880), .A2(net424929), .ZN(net422128) );
  NAND2_X1 U57 ( .A1(net422128), .A2(net424928), .ZN(net425847) );
  AND2_X1 U58 ( .A1(n12), .A2(n11), .ZN(net424929) );
  NOR2_X1 U59 ( .A1(net409390), .A2(n15), .ZN(n12) );
  NAND2_X1 U60 ( .A1(net409394), .A2(net409392), .ZN(n15) );
  AND2_X2 U61 ( .A1(net409418), .A2(net424901), .ZN(net424928) );
  NOR2_X2 U62 ( .A1(n14), .A2(n13), .ZN(net424901) );
  NAND2_X1 U63 ( .A1(net409397), .A2(net409398), .ZN(n13) );
  NAND2_X1 U64 ( .A1(net409400), .A2(net409399), .ZN(n14) );
  INV_X1 U65 ( .A(net409395), .ZN(net409418) );
  OAI21_X1 U66 ( .B1(net412777), .B2(net412829), .A(net409418), .ZN(net412849)
         );
  NAND4_X1 U67 ( .A1(net409419), .A2(net409420), .A3(net409421), .A4(net409422), .ZN(net409395) );
  NAND2_X1 U68 ( .A1(net424880), .A2(net409423), .ZN(net409442) );
  NAND2_X1 U69 ( .A1(net409397), .A2(net409393), .ZN(net409403) );
  NAND2_X1 U70 ( .A1(net409391), .A2(net409400), .ZN(net409416) );
  NAND2_X1 U71 ( .A1(net412849), .A2(net409391), .ZN(net424911) );
  CLKBUF_X1 U72 ( .A(net409390), .Z(net412829) );
  NAND2_X1 U73 ( .A1(net409394), .A2(net409398), .ZN(net409407) );
  AOI21_X1 U74 ( .B1(net412807), .B2(net409394), .A(net424857), .ZN(net409401)
         );
  INV_X1 U75 ( .A(net409392), .ZN(net424868) );
  NAND2_X1 U76 ( .A1(net409392), .A2(net409399), .ZN(net409412) );
  INV_X1 U77 ( .A(net409398), .ZN(net424857) );
  NAND2_X1 U78 ( .A1(net424911), .A2(net409400), .ZN(net424910) );
  OAI211_X1 U79 ( .C1(net424868), .C2(net409400), .A(net424869), .B(net409399), 
        .ZN(net412807) );
  NAND2_X1 U80 ( .A1(net409419), .A2(net409426), .ZN(net409431) );
  NAND2_X1 U81 ( .A1(net422175), .A2(n16), .ZN(net409353) );
  INV_X2 U82 ( .A(A[28]), .ZN(n16) );
  NOR2_X2 U83 ( .A1(n18), .A2(n19), .ZN(n17) );
  AOI21_X1 U84 ( .B1(A[26]), .B2(A[27]), .A(net425779), .ZN(n19) );
  INV_X2 U85 ( .A(net409365), .ZN(n18) );
  NAND2_X1 U86 ( .A1(A[28]), .A2(net425779), .ZN(net409352) );
  AND2_X2 U87 ( .A1(net409364), .A2(net409365), .ZN(net425903) );
  OAI21_X1 U88 ( .B1(A[26]), .B2(net425779), .A(net425858), .ZN(net409375) );
  NOR2_X1 U89 ( .A1(net425779), .A2(A[26]), .ZN(net425889) );
  NAND2_X1 U90 ( .A1(A[26]), .A2(net425779), .ZN(net425858) );
  XNOR2_X1 U91 ( .A(net425779), .B(A[27]), .ZN(net425890) );
  NAND2_X1 U92 ( .A1(A[27]), .A2(net425779), .ZN(net425863) );
  INV_X1 U93 ( .A(net409365), .ZN(net425902) );
  NAND2_X1 U94 ( .A1(net409447), .A2(net425920), .ZN(net424880) );
  NOR2_X1 U95 ( .A1(net409452), .A2(net409453), .ZN(net425920) );
  NAND2_X1 U96 ( .A1(net422175), .A2(n20), .ZN(net409393) );
  INV_X2 U97 ( .A(A[23]), .ZN(n20) );
  NAND2_X1 U98 ( .A1(net422175), .A2(n23), .ZN(net409391) );
  INV_X2 U99 ( .A(A[20]), .ZN(n23) );
  NAND4_X1 U100 ( .A1(net409423), .A2(net409424), .A3(net409425), .A4(
        net409426), .ZN(net409390) );
  NAND2_X1 U101 ( .A1(net409338), .A2(n21), .ZN(net409394) );
  INV_X2 U102 ( .A(A[22]), .ZN(n21) );
  INV_X1 U103 ( .A(B[31]), .ZN(net409338) );
  NAND2_X1 U104 ( .A1(net409338), .A2(n22), .ZN(net409392) );
  INV_X2 U105 ( .A(A[21]), .ZN(n22) );
  AND2_X1 U106 ( .A1(net409447), .A2(net409446), .ZN(net412777) );
  INV_X1 U107 ( .A(net409451), .ZN(net409448) );
  INV_X2 U108 ( .A(net409450), .ZN(net409449) );
  OAI21_X1 U109 ( .B1(net409464), .B2(net409451), .A(net409465), .ZN(net409452) );
  NOR2_X1 U110 ( .A1(net409452), .A2(net409453), .ZN(net409446) );
  INV_X1 U111 ( .A(net409486), .ZN(net409464) );
  CLKBUF_X1 U112 ( .A(net409464), .Z(net412860) );
  OAI211_X1 U113 ( .C1(net409487), .C2(net409488), .A(n24), .B(net409490), 
        .ZN(net409486) );
  NAND2_X1 U114 ( .A1(net422162), .A2(n25), .ZN(n24) );
  OR2_X1 U115 ( .A1(B[11]), .A2(A[11]), .ZN(n25) );
  NAND2_X1 U116 ( .A1(net409494), .A2(net409294), .ZN(net409488) );
  NAND2_X1 U117 ( .A1(net412844), .A2(net409495), .ZN(net409487) );
  NAND2_X1 U118 ( .A1(net409295), .A2(net409298), .ZN(net409495) );
  AOI21_X1 U119 ( .B1(net409454), .B2(net409455), .A(net409456), .ZN(net409453) );
  INV_X1 U120 ( .A(net409457), .ZN(net409456) );
  OAI21_X1 U121 ( .B1(net409458), .B2(net409459), .A(net409460), .ZN(net409454) );
  INV_X2 U122 ( .A(net409461), .ZN(net409459) );
  NOR2_X1 U123 ( .A1(net409462), .A2(net409463), .ZN(net409458) );
  INV_X1 U124 ( .A(net409467), .ZN(net409462) );
  OAI21_X1 U125 ( .B1(net409474), .B2(net409462), .A(net409461), .ZN(net409471) );
  OAI21_X1 U126 ( .B1(net412803), .B2(net409450), .A(net412860), .ZN(net409481) );
  NAND2_X1 U127 ( .A1(net409465), .A2(net409457), .ZN(net409468) );
  NAND2_X1 U128 ( .A1(net409490), .A2(net412844), .ZN(net409498) );
  INV_X4 U129 ( .A(net422162), .ZN(net409493) );
  NAND2_X1 U130 ( .A1(net409457), .A2(n26), .ZN(net409451) );
  AND3_X1 U131 ( .A1(net409467), .A2(net409466), .A3(net409460), .ZN(n26) );
  NAND4_X1 U132 ( .A1(net409494), .A2(net412844), .A3(net422158), .A4(
        net409299), .ZN(net409450) );
  CLKBUF_X1 U133 ( .A(net409294), .Z(net422158) );
  CLKBUF_X1 U134 ( .A(net422158), .Z(net412854) );
  NAND2_X1 U135 ( .A1(net409461), .A2(net409467), .ZN(net409478) );
  INV_X1 U136 ( .A(net409466), .ZN(net409479) );
  NAND2_X1 U137 ( .A1(net409463), .A2(net409466), .ZN(net409484) );
  NAND2_X1 U138 ( .A1(net409460), .A2(net409471), .ZN(net409470) );
  NAND2_X1 U139 ( .A1(net409455), .A2(net409460), .ZN(net409473) );
  INV_X1 U140 ( .A(net409494), .ZN(net409501) );
  NAND2_X1 U141 ( .A1(net409493), .A2(net409494), .ZN(net409505) );
  NAND2_X1 U142 ( .A1(net412837), .A2(net409311), .ZN(net409313) );
  INV_X1 U143 ( .A(B[4]), .ZN(net409531) );
  INV_X1 U144 ( .A(A[4]), .ZN(net409532) );
  NAND2_X1 U145 ( .A1(net412826), .A2(A[4]), .ZN(net409316) );
  NAND2_X2 U146 ( .A1(net409321), .A2(net409322), .ZN(net409317) );
  XNOR2_X1 U147 ( .A(net425779), .B(A[30]), .ZN(net421930) );
  NOR2_X1 U148 ( .A1(net425779), .A2(A[30]), .ZN(net421914) );
  NAND2_X1 U149 ( .A1(net425779), .A2(A[30]), .ZN(net421921) );
  NAND2_X2 U150 ( .A1(n27), .A2(n28), .ZN(net409304) );
  INV_X2 U151 ( .A(A[6]), .ZN(n28) );
  INV_X1 U152 ( .A(B[6]), .ZN(n27) );
  NAND2_X1 U153 ( .A1(B[6]), .A2(A[6]), .ZN(net409303) );
  NAND2_X1 U154 ( .A1(B[5]), .A2(A[5]), .ZN(net409311) );
  OR2_X2 U155 ( .A1(B[5]), .A2(A[5]), .ZN(net409319) );
  OAI21_X1 U156 ( .B1(n33), .B2(net425889), .A(net425858), .ZN(n30) );
  XNOR2_X1 U157 ( .A(n30), .B(net425890), .ZN(SUM[27]) );
  OR2_X1 U158 ( .A1(net425902), .A2(net409363), .ZN(n31) );
  NAND2_X1 U159 ( .A1(net425847), .A2(net425903), .ZN(n32) );
  AND2_X2 U160 ( .A1(n32), .A2(n31), .ZN(n29) );
  AND2_X1 U161 ( .A1(n32), .A2(n34), .ZN(n33) );
  AND2_X1 U162 ( .A1(net409362), .A2(n31), .ZN(n34) );
  NAND2_X1 U163 ( .A1(A[25]), .A2(net425779), .ZN(net409362) );
  NAND2_X1 U164 ( .A1(net422175), .A2(n35), .ZN(net409365) );
  INV_X2 U165 ( .A(A[25]), .ZN(n35) );
  NAND2_X1 U166 ( .A1(net422175), .A2(n36), .ZN(net409364) );
  INV_X2 U167 ( .A(A[24]), .ZN(n36) );
  NAND2_X1 U168 ( .A1(A[24]), .A2(net425779), .ZN(net409363) );
  INV_X2 U169 ( .A(net424910), .ZN(net421184) );
  INV_X1 U170 ( .A(net424932), .ZN(net412845) );
  CLKBUF_X1 U171 ( .A(net412777), .Z(net424932) );
  NAND2_X1 U172 ( .A1(net409470), .A2(net409455), .ZN(net409469) );
  INV_X1 U173 ( .A(net409327), .ZN(n42) );
  AND2_X1 U174 ( .A1(B[10]), .A2(A[10]), .ZN(net422162) );
  INV_X1 U175 ( .A(net409531), .ZN(net422154) );
  CLKBUF_X1 U176 ( .A(net409295), .Z(net422152) );
  CLKBUF_X1 U177 ( .A(net409471), .Z(net422148) );
  OAI21_X1 U178 ( .B1(net409479), .B2(net409480), .A(net409463), .ZN(n37) );
  CLKBUF_X1 U179 ( .A(net409298), .Z(net422142) );
  INV_X1 U180 ( .A(n43), .ZN(n38) );
  XNOR2_X1 U181 ( .A(net409357), .B(net409358), .ZN(SUM[28]) );
  AND2_X1 U182 ( .A1(net409442), .A2(net409422), .ZN(n39) );
  CLKBUF_X1 U183 ( .A(n60), .Z(n40) );
  INV_X1 U184 ( .A(net421184), .ZN(net409410) );
  AOI21_X1 U185 ( .B1(net421916), .B2(net421917), .A(net421914), .ZN(n41) );
  XNOR2_X1 U186 ( .A(n41), .B(n42), .ZN(SUM[31]) );
  INV_X1 U187 ( .A(net421857), .ZN(net412835) );
  CLKBUF_X1 U188 ( .A(net421857), .Z(net409368) );
  CLKBUF_X1 U189 ( .A(net422154), .Z(net412826) );
  XNOR2_X1 U190 ( .A(n65), .B(n63), .ZN(SUM[17]) );
  AND2_X1 U191 ( .A1(net409531), .A2(net409532), .ZN(n43) );
  NAND2_X1 U192 ( .A1(net409316), .A2(n38), .ZN(net409320) );
  INV_X1 U193 ( .A(net409328), .ZN(net409327) );
  XNOR2_X1 U194 ( .A(net425779), .B(A[31]), .ZN(net409328) );
  INV_X1 U195 ( .A(net409480), .ZN(net412863) );
  NAND2_X1 U196 ( .A1(n69), .A2(n70), .ZN(net409460) );
  OAI21_X1 U197 ( .B1(net409479), .B2(net409480), .A(net409463), .ZN(net409475) );
  OR2_X1 U198 ( .A1(B[9]), .A2(A[9]), .ZN(net409294) );
  OR2_X2 U199 ( .A1(B[10]), .A2(A[10]), .ZN(net409494) );
  OR2_X2 U200 ( .A1(B[13]), .A2(A[13]), .ZN(net409467) );
  OR2_X1 U201 ( .A1(B[11]), .A2(A[11]), .ZN(net412844) );
  CLKBUF_X1 U202 ( .A(B[11]), .Z(net412839) );
  OAI21_X1 U203 ( .B1(net409506), .B2(n76), .A(net422152), .ZN(n75) );
  INV_X1 U204 ( .A(net409310), .ZN(net412837) );
  OAI21_X1 U205 ( .B1(A[1]), .B2(B[1]), .A(n52), .ZN(n56) );
  NOR2_X1 U206 ( .A1(A[1]), .A2(B[1]), .ZN(n50) );
  NAND2_X1 U207 ( .A1(B[1]), .A2(A[1]), .ZN(n52) );
  OAI211_X1 U208 ( .C1(n80), .C2(n81), .A(n82), .B(n53), .ZN(net409323) );
  XNOR2_X1 U209 ( .A(net409412), .B(net409410), .ZN(SUM[21]) );
  XNOR2_X1 U210 ( .A(net409468), .B(net409469), .ZN(SUM[15]) );
  NAND2_X1 U211 ( .A1(n59), .A2(net409420), .ZN(n58) );
  NAND2_X1 U212 ( .A1(net409420), .A2(net409425), .ZN(n62) );
  OAI21_X1 U213 ( .B1(n39), .B2(net409438), .A(net409421), .ZN(n60) );
  NAND2_X1 U214 ( .A1(net409421), .A2(net409424), .ZN(n65) );
  NAND2_X1 U215 ( .A1(net409442), .A2(net409422), .ZN(n63) );
  NAND2_X1 U216 ( .A1(net409422), .A2(net409423), .ZN(n67) );
  CLKBUF_X1 U217 ( .A(B[13]), .Z(n44) );
  NAND2_X1 U218 ( .A1(B[12]), .A2(A[12]), .ZN(net409463) );
  INV_X1 U219 ( .A(B[12]), .ZN(n71) );
  NAND2_X1 U220 ( .A1(n44), .A2(A[13]), .ZN(net409461) );
  NAND2_X1 U221 ( .A1(B[14]), .A2(A[14]), .ZN(net409455) );
  INV_X1 U222 ( .A(B[14]), .ZN(n69) );
  NAND2_X1 U223 ( .A1(net422152), .A2(net412854), .ZN(n45) );
  NAND2_X1 U224 ( .A1(B[9]), .A2(A[9]), .ZN(net409295) );
  NAND2_X1 U225 ( .A1(net409531), .A2(net409532), .ZN(net409318) );
  NAND2_X1 U226 ( .A1(net409299), .A2(net422142), .ZN(n47) );
  NAND2_X1 U227 ( .A1(n77), .A2(net422142), .ZN(n46) );
  OAI21_X1 U228 ( .B1(A[2]), .B2(B[2]), .A(n53), .ZN(n48) );
  NAND2_X1 U229 ( .A1(B[2]), .A2(A[2]), .ZN(n53) );
  OAI211_X1 U230 ( .C1(A[2]), .C2(B[2]), .A(A[1]), .B(B[1]), .ZN(n82) );
  OAI22_X1 U231 ( .A1(A[1]), .A2(B[1]), .B1(A[2]), .B2(B[2]), .ZN(n80) );
  NAND2_X1 U232 ( .A1(B[8]), .A2(A[8]), .ZN(net409298) );
  INV_X1 U233 ( .A(B[8]), .ZN(n78) );
  CLKBUF_X1 U234 ( .A(net412849), .Z(net412813) );
  XNOR2_X1 U235 ( .A(net409407), .B(net412807), .ZN(SUM[22]) );
  OR2_X1 U236 ( .A1(B[31]), .A2(A[15]), .ZN(net409457) );
  NAND2_X1 U237 ( .A1(net412839), .A2(A[11]), .ZN(net409490) );
  XNOR2_X1 U238 ( .A(net409431), .B(n58), .ZN(SUM[19]) );
  XNOR2_X1 U239 ( .A(n62), .B(n40), .ZN(SUM[18]) );
  NAND2_X1 U240 ( .A1(net409425), .A2(n60), .ZN(n59) );
  XNOR2_X1 U241 ( .A(net409478), .B(n37), .ZN(SUM[13]) );
  NAND2_X1 U242 ( .A1(n71), .A2(n72), .ZN(net409466) );
  NAND2_X1 U243 ( .A1(net409382), .A2(net409363), .ZN(n54) );
  INV_X1 U244 ( .A(net412803), .ZN(net412778) );
  XNOR2_X1 U245 ( .A(net409401), .B(net409402), .ZN(SUM[23]) );
  XNOR2_X1 U246 ( .A(net409416), .B(net412813), .ZN(SUM[20]) );
  XNOR2_X1 U247 ( .A(net412793), .B(net409346), .ZN(SUM[29]) );
  XNOR2_X1 U248 ( .A(net409368), .B(net409383), .ZN(SUM[24]) );
  XNOR2_X1 U249 ( .A(n47), .B(net412778), .ZN(SUM[8]) );
  NAND2_X1 U250 ( .A1(net412841), .A2(net409299), .ZN(n77) );
  XNOR2_X1 U251 ( .A(n54), .B(net409380), .ZN(SUM[25]) );
  XNOR2_X1 U252 ( .A(net412845), .B(n67), .ZN(SUM[16]) );
  XNOR2_X1 U253 ( .A(net422133), .B(net409375), .ZN(SUM[26]) );
  NAND2_X1 U254 ( .A1(A[23]), .A2(net425779), .ZN(net409397) );
  NAND2_X1 U255 ( .A1(A[19]), .A2(net425779), .ZN(net409419) );
  NAND2_X1 U256 ( .A1(A[22]), .A2(B[31]), .ZN(net409398) );
  NAND2_X1 U257 ( .A1(A[21]), .A2(net425779), .ZN(net409399) );
  NAND2_X1 U258 ( .A1(A[18]), .A2(B[31]), .ZN(net409420) );
  NAND2_X1 U259 ( .A1(A[20]), .A2(B[31]), .ZN(net409400) );
  NAND2_X1 U260 ( .A1(A[17]), .A2(B[31]), .ZN(net409421) );
  NAND2_X1 U261 ( .A1(A[16]), .A2(B[31]), .ZN(net409422) );
  NAND2_X1 U262 ( .A1(net409338), .A2(n68), .ZN(net409423) );
  NAND2_X1 U263 ( .A1(net409338), .A2(n61), .ZN(net409426) );
  NAND2_X1 U264 ( .A1(net409338), .A2(n66), .ZN(net409424) );
  NAND2_X1 U265 ( .A1(net409338), .A2(n64), .ZN(net409425) );
  NAND2_X1 U266 ( .A1(A[15]), .A2(B[31]), .ZN(net409465) );
  XNOR2_X2 U267 ( .A(n45), .B(n46), .ZN(SUM[9]) );
  XNOR2_X2 U268 ( .A(net409300), .B(net409301), .ZN(SUM[7]) );
  NAND2_X2 U269 ( .A1(net409304), .A2(net409305), .ZN(net409302) );
  XNOR2_X2 U270 ( .A(net409308), .B(net409305), .ZN(SUM[6]) );
  INV_X1 U271 ( .A(net409312), .ZN(net409309) );
  XNOR2_X2 U272 ( .A(net409313), .B(net409312), .ZN(SUM[5]) );
  OAI21_X2 U273 ( .B1(n43), .B2(net409315), .A(net409316), .ZN(net409312) );
  INV_X1 U274 ( .A(net409317), .ZN(net409315) );
  XNOR2_X2 U275 ( .A(net409320), .B(net409317), .ZN(SUM[4]) );
  XNOR2_X1 U276 ( .A(net409325), .B(net412864), .ZN(SUM[3]) );
  XNOR2_X1 U277 ( .A(n48), .B(n49), .ZN(SUM[2]) );
  OAI21_X2 U278 ( .B1(n50), .B2(n51), .A(n52), .ZN(n49) );
  NAND2_X1 U279 ( .A1(A[0]), .A2(B[0]), .ZN(n51) );
  INV_X1 U280 ( .A(net409403), .ZN(net409402) );
  XNOR2_X1 U281 ( .A(n55), .B(n56), .ZN(SUM[1]) );
  INV_X1 U282 ( .A(n57), .ZN(n55) );
  INV_X2 U283 ( .A(A[19]), .ZN(n61) );
  INV_X1 U284 ( .A(net409424), .ZN(net409438) );
  INV_X2 U285 ( .A(A[18]), .ZN(n64) );
  INV_X2 U286 ( .A(A[17]), .ZN(n66) );
  INV_X2 U287 ( .A(A[16]), .ZN(n68) );
  XNOR2_X1 U288 ( .A(net422148), .B(net409473), .ZN(SUM[14]) );
  INV_X1 U289 ( .A(net409475), .ZN(net409474) );
  INV_X2 U290 ( .A(A[14]), .ZN(n70) );
  INV_X1 U291 ( .A(net409481), .ZN(net409480) );
  XNOR2_X1 U292 ( .A(net409484), .B(net412863), .ZN(SUM[12]) );
  INV_X2 U293 ( .A(A[12]), .ZN(n72) );
  XNOR2_X1 U294 ( .A(net409498), .B(n73), .ZN(SUM[11]) );
  OAI21_X1 U295 ( .B1(n74), .B2(net409501), .A(net409493), .ZN(n73) );
  INV_X1 U296 ( .A(n75), .ZN(n74) );
  XNOR2_X2 U297 ( .A(net409505), .B(n75), .ZN(SUM[10]) );
  INV_X1 U298 ( .A(n46), .ZN(n76) );
  NAND2_X2 U299 ( .A1(n78), .A2(n79), .ZN(net409299) );
  INV_X2 U300 ( .A(A[8]), .ZN(n79) );
  NAND2_X2 U301 ( .A1(B[3]), .A2(A[3]), .ZN(net409322) );
  NAND2_X1 U302 ( .A1(B[0]), .A2(A[0]), .ZN(n81) );
  NAND2_X2 U303 ( .A1(n83), .A2(n84), .ZN(net409324) );
  INV_X2 U304 ( .A(A[3]), .ZN(n84) );
  INV_X2 U305 ( .A(B[3]), .ZN(n83) );
  INV_X1 U306 ( .A(net412854), .ZN(net409506) );
  INV_X2 U307 ( .A(n85), .ZN(SUM[0]) );
  OAI21_X2 U308 ( .B1(A[0]), .B2(B[0]), .A(n57), .ZN(n85) );
  NAND2_X2 U309 ( .A1(B[0]), .A2(A[0]), .ZN(n57) );
endmodule


module carry_sel_bk_NB4_48 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U12 ( .A(n30), .ZN(n5) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
endmodule


module carry_sel_bk_NB4_31 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n7) );
  INV_X1 U2 ( .A(n12), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI22_X1 U4 ( .A1(n9), .A2(n1), .B1(Ci), .B2(n8), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n10), .A2(n7), .B1(n5), .B2(n4), .ZN(n9) );
  AOI22_X1 U6 ( .A1(n7), .A2(n30), .B1(n6), .B2(n5), .ZN(n8) );
  NAND2_X1 U7 ( .A1(n3), .A2(n13), .ZN(n5) );
  OAI22_X1 U8 ( .A1(n36), .A2(n1), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(n37), .A2(n34), .B1(n33), .B2(n12), .ZN(n36) );
  AOI22_X1 U10 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U11 ( .A1(n11), .A2(n39), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n1), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U16 ( .A(Ci), .B(n2), .ZN(S[0]) );
  NAND2_X1 U17 ( .A1(n4), .A2(n30), .ZN(n2) );
  OAI21_X1 U18 ( .B1(n31), .B2(n30), .A(n13), .ZN(n32) );
  OAI21_X1 U19 ( .B1(n10), .B2(n31), .A(n13), .ZN(n12) );
  OAI21_X1 U20 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U21 ( .A(n10), .ZN(n4) );
  INV_X1 U22 ( .A(n30), .ZN(n6) );
  INV_X1 U23 ( .A(n40), .ZN(n11) );
  INV_X1 U24 ( .A(n31), .ZN(n3) );
  NOR2_X1 U25 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U27 ( .A1(B[0]), .A2(A[0]), .ZN(n10) );
  NAND2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U29 ( .A1(B[1]), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  INV_X1 U31 ( .A(Ci), .ZN(n1) );
endmodule


module carry_sel_bk_NB4_32 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U12 ( .A(n30), .ZN(n5) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_24 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U12 ( .A(n30), .ZN(n5) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_16 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U12 ( .A(n30), .ZN(n5) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_33 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_25 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_22 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_14 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_57 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
endmodule


module carry_sel_bk_NB4_56 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
endmodule


module carry_sel_bk_NB4_13 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
endmodule


module carry_sel_bk_NB4_60 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_53 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_52 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_45 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_44 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_43 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_37 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_36 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_35 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_28 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_27 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_20 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_19 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_54 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_30 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_26 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_18 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI21_X1 U5 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  AOI22_X1 U8 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U9 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  INV_X1 U11 ( .A(n30), .ZN(n5) );
  XNOR2_X1 U12 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U13 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NAND2_X1 U16 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U17 ( .A(n31), .ZN(n2) );
  NAND2_X1 U18 ( .A1(n10), .A2(n39), .ZN(n33) );
  INV_X1 U19 ( .A(n40), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U21 ( .A(n9), .ZN(n3) );
  NOR2_X1 U22 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U23 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U24 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U25 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U27 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  XNOR2_X1 U28 ( .A(Ci), .B(n1), .ZN(S[0]) );
  OAI22_X1 U29 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  OAI22_X1 U30 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  OAI22_X1 U31 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
endmodule


module carry_sel_bk_NB4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI21_X1 U5 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  AOI22_X1 U8 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  INV_X1 U9 ( .A(n30), .ZN(n5) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  XNOR2_X1 U12 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U13 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NAND2_X1 U16 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U17 ( .A(n31), .ZN(n2) );
  NAND2_X1 U18 ( .A1(n10), .A2(n39), .ZN(n33) );
  INV_X1 U19 ( .A(n40), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U21 ( .A(n9), .ZN(n3) );
  NOR2_X1 U22 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U23 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U24 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U27 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  XNOR2_X1 U28 ( .A(Ci), .B(n1), .ZN(S[0]) );
  OAI22_X1 U29 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  OAI22_X1 U30 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  OAI22_X1 U31 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
endmodule


module G_78 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2, n1;

  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n1) );
  INV_X1 U3 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Gij) );
endmodule


module G_71 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_70 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_69 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_68 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_67 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_66 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_65 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_64 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_63 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_62 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_61 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_60 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_59 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_58 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_57 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_56 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_55 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_54 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_53 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_52 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_51 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_50 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_49 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_48 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_47 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_46 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_45 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_44 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_43 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_42 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_41 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_40 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_39 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_38 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_37 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_36 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_35 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_34 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_33 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_32 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_31 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_30 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_29 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_28 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_27 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_26 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_25 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_24 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_23 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_22 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_21 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_20 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_19 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_18 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_17 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_16 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_15 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_14 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_13 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_12 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_11 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_10 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_9 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_8 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_7 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_6 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_5 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_4 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_3 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_2 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_1 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module G_0 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module blockPG_230 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  OR2_X1 U2 ( .A1(Gik), .A2(n2), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
endmodule


module blockPG_227 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_226 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_240 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module blockPG_236 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module blockPG_225 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module blockPG_219 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  NAND2_X1 U1 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_235 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_234 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_231 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_224 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_223 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_222 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_216 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_47 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_228 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_221 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_215 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_214 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_213 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_212 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_211 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_209 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_208 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_207 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_204 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_203 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_199 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_198 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_197 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_196 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_195 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_194 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_192 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_188 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_187 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_186 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_185 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_184 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_182 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_181 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_180 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_177 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_176 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_172 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_171 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_170 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_169 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_168 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_167 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_165 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_161 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_160 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_159 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_158 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_157 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_155 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_154 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_153 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_150 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_149 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_145 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_144 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_143 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_142 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_141 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_140 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_138 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_134 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_133 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_132 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_131 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_130 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_128 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_127 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_126 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_123 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_122 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_118 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_117 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_116 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_115 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_114 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_113 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_111 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_107 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_106 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_105 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_104 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_101 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_100 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_99 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_96 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_95 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_91 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_90 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_89 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_88 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_87 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_86 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_84 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_80 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_79 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_78 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_77 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_76 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_74 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_73 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_72 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_69 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_68 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_64 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_63 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_62 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_61 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_60 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_59 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_57 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_53 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_52 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_51 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_50 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_49 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_46 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_45 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_42 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_41 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_37 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_36 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_35 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_34 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_33 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_32 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_30 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_26 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_25 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_24 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_23 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_22 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_19 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_18 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_15 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_14 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_10 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_9 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_8 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_7 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_6 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_5 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_3 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_210 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_206 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_205 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_202 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_201 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_191 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_183 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_179 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_178 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_175 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_174 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_164 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_156 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_152 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_151 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_148 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_147 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_137 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_129 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_125 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_124 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_121 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_120 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_110 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_102 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_98 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_97 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_94 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_93 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_83 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_75 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_71 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_70 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_67 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_66 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_56 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_48 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_44 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_43 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_40 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_39 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_29 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_20 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_17 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_16 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_13 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_12 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_2 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_200 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_193 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_190 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_189 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_173 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_166 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_163 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_162 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_146 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_139 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_136 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_135 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_119 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_112 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_109 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_108 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_92 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_85 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_82 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_81 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_65 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_58 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_55 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_54 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_38 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_31 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_28 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_27 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_21 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_11 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_4 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_1 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_0 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module pg_net_285 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module pg_net_275 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_274 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_278 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module pg_net_270 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module pg_net_262 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module pg_net_281 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p) );
endmodule


module pg_net_277 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p) );
endmodule


module pg_net_273 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p) );
endmodule


module pg_net_269 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p) );
endmodule


module pg_net_265 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p) );
endmodule


module pg_net_261 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p) );
endmodule


module pg_net_279 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_276 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(n2), .ZN(g) );
  CLKBUF_X1 U3 ( .A(b), .Z(n2) );
endmodule


module pg_net_272 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_271 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_268 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_267 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_266 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_264 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_263 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_260 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_258 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_257 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_256 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_255 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_254 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_253 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_252 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_251 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_250 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_249 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_248 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_247 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_246 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_245 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_244 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_243 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_242 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_241 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_240 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_239 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_238 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_237 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_236 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_235 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_234 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_233 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_232 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_231 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_230 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_229 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_228 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_227 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_226 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_225 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_224 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_223 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_222 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_221 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_220 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_219 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_218 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_217 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_216 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_215 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_214 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_213 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_212 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_211 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_210 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_209 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_208 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_207 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_206 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_205 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_204 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_203 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_202 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_201 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_200 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_199 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_198 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_197 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_196 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_195 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_194 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_193 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_192 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_191 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_190 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_189 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_188 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_187 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_186 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_185 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_184 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_183 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_182 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_181 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_180 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_179 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_178 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_177 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_176 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_175 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_174 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_173 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_172 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_171 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_170 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_169 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_168 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_167 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_166 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_165 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_164 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_163 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_162 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_161 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_160 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_159 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_158 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_157 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_156 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_155 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_154 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_153 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_152 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_151 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_150 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_149 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_148 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_147 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_146 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_145 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_144 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_143 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_142 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_141 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_140 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_139 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_138 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_137 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_136 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_135 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_134 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_133 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_132 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_131 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_130 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_129 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_128 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_127 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_126 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_125 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_124 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_123 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_122 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_121 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_120 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_119 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_118 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_117 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_116 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_115 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_114 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_113 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_112 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_111 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_110 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_109 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_108 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_107 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_106 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_105 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_104 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_103 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_102 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_101 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_100 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_99 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_98 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_97 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_96 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_95 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_94 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_93 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_92 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_91 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_90 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_89 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_88 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_87 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_86 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_85 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_84 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_83 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_82 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_81 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_80 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_79 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_78 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_77 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_76 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_75 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_74 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_73 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_72 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_71 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_70 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_69 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_68 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_67 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_66 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_65 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_64 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_63 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_62 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_61 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_60 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_59 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_58 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_57 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_56 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_55 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_54 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_53 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_52 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_51 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_50 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_49 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_48 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_47 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_46 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_45 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_44 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_43 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_42 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_41 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_40 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_39 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_38 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_37 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_36 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_35 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_34 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_33 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_32 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_31 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_30 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_28 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_27 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_26 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_25 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_24 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_23 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_22 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_21 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_20 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_19 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_18 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_17 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_15 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_14 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_13 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_12 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_11 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_10 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_9 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_8 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_7 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_6 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_5 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_0 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module CSTgen_CW4_NB32_6 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_223 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_222 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_221 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_220 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_219 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_218 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_217 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_216 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_215 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_214 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_213 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_212 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_211 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_210 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_209 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_208 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_207 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_206 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_205 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_204 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_203 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_202 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_201 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_200 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_199 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_198 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_197 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_196 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_195 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_194 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_193 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_192 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_188 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_62 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_187 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_186 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_185 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_184 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_183 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_182 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_181 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_180 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_179 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_178 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_177 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_176 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_175 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_174 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_61 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_173 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_172 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_171 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_170 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_169 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_168 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_167 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_60 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_166 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_165 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_164 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_59 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_58 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_163 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_162 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_57 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_56 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_55 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_54 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module CSTgen_CW4_NB32_5 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_191 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_190 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_189 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_188 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_187 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_186 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_185 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_184 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_183 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_182 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_181 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_180 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_179 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_178 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_177 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_176 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_175 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_174 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_173 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_172 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_171 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_170 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_169 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_168 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_167 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_166 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_165 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_164 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_163 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_162 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_161 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_160 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_161 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_53 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_160 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_159 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_158 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_157 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_156 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_155 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_154 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_153 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_152 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_151 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_150 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_149 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_148 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_147 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_52 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_146 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_145 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_144 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_143 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_142 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_141 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_140 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_51 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_139 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_138 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_137 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_50 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_49 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_136 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_135 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_48 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_47 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_46 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_45 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module CSTgen_CW4_NB32_4 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_159 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_158 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_157 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_156 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_155 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_154 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_153 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_152 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_151 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_150 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_149 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_148 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_147 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_146 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_145 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_144 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_143 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_142 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_141 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_140 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_139 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_138 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_137 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_136 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_135 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_134 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_133 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_132 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_131 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_130 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_129 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_128 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_134 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_44 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_133 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_132 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_131 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_130 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_129 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_128 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_127 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_126 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_125 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_124 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_123 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_122 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_121 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_120 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_43 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_119 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_118 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_117 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_116 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_115 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_114 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_113 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_42 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_112 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_111 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_110 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_41 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_40 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_109 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_108 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_39 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_38 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_37 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_36 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module CSTgen_CW4_NB32_2 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_95 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_94 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_93 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_92 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_91 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_90 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_89 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_88 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_87 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_86 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_85 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_84 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_83 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_82 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_81 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_80 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_79 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_78 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_77 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_76 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_75 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_74 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_73 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_72 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_71 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_70 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_69 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_68 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_67 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_66 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_65 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_64 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_80 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_26 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_79 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_78 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_77 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_76 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_75 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_74 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_73 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_72 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_71 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_70 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_69 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_68 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_67 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_66 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_25 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_65 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_64 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_63 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_62 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_61 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_60 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_59 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_24 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_58 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_57 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_56 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_23 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_22 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_55 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_54 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_21 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_20 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_19 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_18 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module MUX21_generic_NB32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  CLKBUF_X1 U1 ( .A(SEL), .Z(n3) );
  CLKBUF_X3 U2 ( .A(SEL), .Z(n1) );
  CLKBUF_X3 U3 ( .A(SEL), .Z(n2) );
  MUX2_X1 U4 ( .A(B[0]), .B(A[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(B[1]), .B(A[1]), .S(n1), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(B[2]), .B(A[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U7 ( .A(B[3]), .B(A[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U8 ( .A(B[4]), .B(A[4]), .S(n1), .Z(Y[4]) );
  MUX2_X1 U9 ( .A(B[5]), .B(A[5]), .S(n1), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(B[6]), .B(A[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(B[7]), .B(A[7]), .S(n1), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(B[8]), .B(A[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(B[9]), .B(A[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(B[10]), .B(A[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(B[11]), .B(A[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(B[12]), .B(A[12]), .S(n2), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(B[13]), .B(A[13]), .S(n2), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(B[14]), .B(A[14]), .S(n2), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(B[15]), .B(A[15]), .S(n2), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(B[16]), .B(A[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(B[17]), .B(A[17]), .S(n2), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(B[18]), .B(A[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(B[19]), .B(A[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(B[20]), .B(A[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(B[21]), .B(A[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(B[22]), .B(A[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(B[23]), .B(A[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(B[24]), .B(A[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(B[25]), .B(A[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(B[26]), .B(A[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(B[27]), .B(A[27]), .S(n3), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(B[28]), .B(A[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(B[29]), .B(A[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(B[30]), .B(A[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(B[31]), .B(A[31]), .S(n3), .Z(Y[31]) );
endmodule


module FD_NB32_2 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n33, n34, n35;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n35), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n35), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n34), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n34), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n34), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n34), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n33), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n33), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n33), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n33), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n33), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n33), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n33), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n33), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n33), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n33), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n33), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n33), .Q(Q[0]) );
  BUF_X1 U3 ( .A(RESET), .Z(n33) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
endmodule


module FD_NB32_1 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n33, n34, n35;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n35), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n35), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n34), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n34), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n34), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n34), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n33), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n33), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n33), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n33), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n33), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n33), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n33), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n33), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n33), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n33), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n33), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n33), .Q(Q[0]) );
  BUF_X1 U3 ( .A(RESET), .Z(n33) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
endmodule


module FD_NB32_0 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n33, n34, n35;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n35), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n35), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n34), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n34), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n34), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n34), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n33), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n33), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n33), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n33), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n33), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n33), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n33), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n33), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n33), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n33), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n33), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n33), .Q(Q[0]) );
  BUF_X1 U3 ( .A(RESET), .Z(n33) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
endmodule


module FD_INJ_NB1_0 ( CK, RESET, INJ_ZERO, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   \TMP_D[0] ;

  DFFR_X1 \Q_reg[0]  ( .D(\TMP_D[0] ), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[0]), .ZN(\TMP_D[0] ) );
endmodule


module FD_NB2_1 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB2_0 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_20 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_19 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_18 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_17 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_16 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_15 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_14 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_13 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_12 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_11 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_10 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_9 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_8 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_7 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_6 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_5 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_4 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_3 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_2 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_1 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_0 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_1 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_0 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module carry_sel_bk_NB4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI21_X1 U5 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI22_X1 U7 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U8 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U9 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U10 ( .A1(n10), .A2(n39), .ZN(n33) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  INV_X1 U12 ( .A(n30), .ZN(n5) );
  AOI22_X1 U13 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U16 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U17 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NAND2_X1 U18 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U19 ( .A(n31), .ZN(n2) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U21 ( .A(n9), .ZN(n3) );
  INV_X1 U22 ( .A(n40), .ZN(n10) );
  NOR2_X1 U23 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U24 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U28 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  XNOR2_X1 U29 ( .A(Ci), .B(n1), .ZN(S[0]) );
  OAI22_X1 U30 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  OAI22_X1 U31 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
endmodule


module carry_sel_bk_NB4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI21_X1 U5 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  AOI22_X1 U8 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  INV_X1 U9 ( .A(n30), .ZN(n5) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  XNOR2_X1 U12 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U13 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NAND2_X1 U16 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U17 ( .A(n31), .ZN(n2) );
  NAND2_X1 U18 ( .A1(n10), .A2(n39), .ZN(n33) );
  INV_X1 U19 ( .A(n40), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U21 ( .A(n9), .ZN(n3) );
  NOR2_X1 U22 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U23 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U24 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U27 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  XNOR2_X1 U28 ( .A(Ci), .B(n1), .ZN(S[0]) );
  OAI22_X1 U29 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  OAI22_X1 U30 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  OAI22_X1 U31 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
endmodule


module carry_sel_bk_NB4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI21_X1 U5 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  AOI22_X1 U8 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  INV_X1 U9 ( .A(n30), .ZN(n5) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  XNOR2_X1 U12 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U13 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NAND2_X1 U16 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U17 ( .A(n31), .ZN(n2) );
  NAND2_X1 U18 ( .A1(n10), .A2(n39), .ZN(n33) );
  INV_X1 U19 ( .A(n40), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U21 ( .A(n9), .ZN(n3) );
  NOR2_X1 U22 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U23 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U24 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U27 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  XNOR2_X1 U28 ( .A(Ci), .B(n1), .ZN(S[0]) );
  OAI22_X1 U29 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  OAI22_X1 U30 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  OAI22_X1 U31 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
endmodule


module carry_sel_bk_NB4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI21_X1 U5 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U8 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  AOI22_X1 U9 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  INV_X1 U10 ( .A(n30), .ZN(n5) );
  AOI22_X1 U11 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U13 ( .A(n31), .ZN(n2) );
  NAND2_X1 U14 ( .A1(n10), .A2(n39), .ZN(n33) );
  INV_X1 U15 ( .A(n40), .ZN(n10) );
  NAND2_X1 U16 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U17 ( .A(n9), .ZN(n3) );
  NOR2_X1 U18 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U19 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NAND2_X1 U20 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U22 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U23 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  XNOR2_X1 U24 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U25 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U26 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U27 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U28 ( .A(Ci), .B(n1), .ZN(S[0]) );
  OAI22_X1 U29 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  OAI22_X1 U30 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  OAI22_X1 U31 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
endmodule


module carry_sel_bk_NB4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI21_X1 U5 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U6 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  AOI22_X1 U8 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U9 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  INV_X1 U11 ( .A(n30), .ZN(n5) );
  XNOR2_X1 U12 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U13 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NAND2_X1 U16 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U17 ( .A(n31), .ZN(n2) );
  NAND2_X1 U18 ( .A1(n10), .A2(n39), .ZN(n33) );
  INV_X1 U19 ( .A(n40), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U21 ( .A(n9), .ZN(n3) );
  NOR2_X1 U22 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U23 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U24 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U25 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U27 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  XNOR2_X1 U28 ( .A(Ci), .B(n1), .ZN(S[0]) );
  OAI22_X1 U29 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  OAI22_X1 U30 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  OAI22_X1 U31 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
endmodule


module carry_sel_bk_NB4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n7) );
  INV_X1 U2 ( .A(n12), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI21_X1 U4 ( .B1(n31), .B2(n30), .A(n13), .ZN(n32) );
  OAI21_X1 U5 ( .B1(n10), .B2(n31), .A(n13), .ZN(n12) );
  AOI22_X1 U6 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  AOI22_X1 U7 ( .A1(n37), .A2(n34), .B1(n33), .B2(n12), .ZN(n36) );
  AOI22_X1 U8 ( .A1(n10), .A2(n7), .B1(n5), .B2(n4), .ZN(n9) );
  AOI22_X1 U9 ( .A1(n7), .A2(n30), .B1(n6), .B2(n5), .ZN(n8) );
  INV_X1 U10 ( .A(n30), .ZN(n6) );
  XNOR2_X1 U11 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U12 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  OAI21_X1 U14 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NAND2_X1 U15 ( .A1(n3), .A2(n13), .ZN(n5) );
  INV_X1 U16 ( .A(n31), .ZN(n3) );
  NAND2_X1 U17 ( .A1(n11), .A2(n39), .ZN(n33) );
  INV_X1 U18 ( .A(n40), .ZN(n11) );
  NAND2_X1 U19 ( .A1(n4), .A2(n30), .ZN(n2) );
  INV_X1 U20 ( .A(n10), .ZN(n4) );
  NOR2_X1 U21 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U22 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U23 ( .A1(B[1]), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U24 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n10) );
  NAND2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n9), .A2(n1), .B1(Ci), .B2(n8), .ZN(S[1]) );
  OAI22_X1 U28 ( .A1(n36), .A2(n1), .B1(Ci), .B2(n35), .ZN(S[2]) );
  OAI22_X1 U29 ( .A1(n1), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U30 ( .A(Ci), .B(n2), .ZN(S[0]) );
  INV_X1 U31 ( .A(Ci), .ZN(n1) );
endmodule


module carry_sel_bk_NB4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  XNOR2_X1 U9 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U10 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U11 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U12 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  INV_X1 U13 ( .A(n9), .ZN(n3) );
  INV_X1 U14 ( .A(n30), .ZN(n5) );
  INV_X1 U15 ( .A(n31), .ZN(n2) );
  OAI22_X1 U16 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U17 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U18 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U19 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U20 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U21 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U22 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U23 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NOR2_X1 U24 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  OAI21_X1 U28 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U29 ( .A(n40), .ZN(n10) );
  NOR2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_15 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n7) );
  INV_X1 U2 ( .A(n12), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI22_X1 U4 ( .A1(n9), .A2(n1), .B1(Ci), .B2(n8), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n7), .A2(n30), .B1(n6), .B2(n5), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n10), .A2(n7), .B1(n5), .B2(n4), .ZN(n9) );
  INV_X1 U7 ( .A(n30), .ZN(n6) );
  OAI22_X1 U8 ( .A1(n36), .A2(n1), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(n37), .A2(n34), .B1(n33), .B2(n12), .ZN(n36) );
  AOI22_X1 U10 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U11 ( .A1(n11), .A2(n39), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n1), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U16 ( .A(Ci), .B(n2), .ZN(S[0]) );
  NAND2_X1 U17 ( .A1(n4), .A2(n30), .ZN(n2) );
  OAI21_X1 U18 ( .B1(n31), .B2(n30), .A(n13), .ZN(n32) );
  OAI21_X1 U19 ( .B1(n10), .B2(n31), .A(n13), .ZN(n12) );
  OAI21_X1 U20 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U21 ( .A1(n3), .A2(n13), .ZN(n5) );
  INV_X1 U22 ( .A(n31), .ZN(n3) );
  INV_X1 U23 ( .A(n10), .ZN(n4) );
  INV_X1 U24 ( .A(n40), .ZN(n11) );
  NOR2_X1 U25 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U28 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n10) );
  NAND2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  INV_X1 U31 ( .A(Ci), .ZN(n1) );
endmodule


module carry_sel_bk_NB4_17 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n40), .ZN(n10) );
  INV_X1 U24 ( .A(n30), .ZN(n5) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_21 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  INV_X1 U4 ( .A(n11), .ZN(n37) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U20 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NAND2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NOR2_X1 U27 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NOR2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U29 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NOR2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_23 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n7) );
  INV_X1 U2 ( .A(n32), .ZN(n41) );
  INV_X1 U3 ( .A(n12), .ZN(n37) );
  OAI22_X1 U4 ( .A1(n9), .A2(n1), .B1(Ci), .B2(n8), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n7), .A2(n30), .B1(n6), .B2(n5), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n10), .A2(n7), .B1(n5), .B2(n4), .ZN(n9) );
  INV_X1 U7 ( .A(n30), .ZN(n6) );
  OAI22_X1 U8 ( .A1(n36), .A2(n1), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(n37), .A2(n34), .B1(n33), .B2(n12), .ZN(n36) );
  AOI22_X1 U10 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U11 ( .A1(n11), .A2(n39), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n1), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U16 ( .A(Ci), .B(n2), .ZN(S[0]) );
  NAND2_X1 U17 ( .A1(n4), .A2(n30), .ZN(n2) );
  OAI21_X1 U18 ( .B1(n10), .B2(n31), .A(n13), .ZN(n12) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n13), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U21 ( .A1(n3), .A2(n13), .ZN(n5) );
  INV_X1 U22 ( .A(n31), .ZN(n3) );
  INV_X1 U23 ( .A(n10), .ZN(n4) );
  INV_X1 U24 ( .A(n40), .ZN(n11) );
  NAND2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NOR2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n10) );
  NOR2_X1 U27 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U29 ( .A1(B[1]), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  INV_X1 U31 ( .A(Ci), .ZN(n1) );
endmodule


module carry_sel_bk_NB4_29 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(n11), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI22_X1 U4 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n2), .A2(n12), .ZN(n4) );
  XNOR2_X1 U8 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U9 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U10 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U11 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  INV_X1 U12 ( .A(Ci), .ZN(n46) );
  INV_X1 U13 ( .A(n9), .ZN(n3) );
  INV_X1 U14 ( .A(n30), .ZN(n5) );
  INV_X1 U15 ( .A(n31), .ZN(n2) );
  OAI22_X1 U16 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U17 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U18 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U19 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U20 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U21 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U22 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U23 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  NOR2_X1 U24 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  OAI21_X1 U28 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U29 ( .A(n40), .ZN(n10) );
  NOR2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module blockPG_103 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module carry_sel_bk_NB4_34 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  OAI22_X1 U2 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U3 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U4 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U5 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U6 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U7 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U8 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U9 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  OAI21_X1 U10 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U11 ( .A(Ci), .ZN(n46) );
  INV_X1 U12 ( .A(n11), .ZN(n37) );
  INV_X1 U13 ( .A(n32), .ZN(n41) );
  INV_X1 U14 ( .A(n40), .ZN(n10) );
  OAI22_X1 U15 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U16 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U17 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U18 ( .A1(n2), .A2(n12), .ZN(n4) );
  NOR2_X1 U19 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  XNOR2_X1 U20 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U21 ( .A1(n3), .A2(n30), .ZN(n1) );
  NAND2_X1 U22 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  OAI21_X1 U23 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U24 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  INV_X1 U25 ( .A(n9), .ZN(n3) );
  INV_X1 U26 ( .A(n30), .ZN(n5) );
  INV_X1 U27 ( .A(n31), .ZN(n2) );
  NOR2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_38 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  OAI22_X1 U2 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U3 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U4 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U5 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U6 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U7 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U8 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U9 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  OAI21_X1 U10 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U11 ( .A(Ci), .ZN(n46) );
  INV_X1 U12 ( .A(n11), .ZN(n37) );
  INV_X1 U13 ( .A(n32), .ZN(n41) );
  INV_X1 U14 ( .A(n40), .ZN(n10) );
  OAI22_X1 U15 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U16 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U17 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U18 ( .A1(n2), .A2(n12), .ZN(n4) );
  XNOR2_X1 U19 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  NOR2_X1 U21 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  OAI21_X1 U22 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U23 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  NAND2_X1 U24 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  INV_X1 U25 ( .A(n9), .ZN(n3) );
  INV_X1 U26 ( .A(n30), .ZN(n5) );
  INV_X1 U27 ( .A(n31), .ZN(n2) );
  NOR2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_39 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n7) );
  INV_X1 U2 ( .A(n12), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI22_X1 U4 ( .A1(n9), .A2(n1), .B1(Ci), .B2(n8), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n10), .A2(n7), .B1(n5), .B2(n4), .ZN(n9) );
  AOI22_X1 U6 ( .A1(n7), .A2(n30), .B1(n6), .B2(n5), .ZN(n8) );
  NAND2_X1 U7 ( .A1(n3), .A2(n13), .ZN(n5) );
  OAI22_X1 U8 ( .A1(n36), .A2(n1), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(n37), .A2(n34), .B1(n33), .B2(n12), .ZN(n36) );
  AOI22_X1 U10 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U11 ( .A1(n11), .A2(n39), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n1), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U16 ( .A(Ci), .B(n2), .ZN(S[0]) );
  NAND2_X1 U17 ( .A1(n4), .A2(n30), .ZN(n2) );
  OAI21_X1 U18 ( .B1(n31), .B2(n30), .A(n13), .ZN(n32) );
  OAI21_X1 U19 ( .B1(n10), .B2(n31), .A(n13), .ZN(n12) );
  OAI21_X1 U20 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U21 ( .A(n10), .ZN(n4) );
  INV_X1 U22 ( .A(n30), .ZN(n6) );
  INV_X1 U23 ( .A(n40), .ZN(n11) );
  INV_X1 U24 ( .A(n31), .ZN(n3) );
  NOR2_X1 U25 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U27 ( .A1(B[0]), .A2(A[0]), .ZN(n10) );
  NAND2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U29 ( .A1(B[1]), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  INV_X1 U31 ( .A(Ci), .ZN(n1) );
endmodule


module carry_sel_bk_NB4_40 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_41 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_42 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U12 ( .A(n30), .ZN(n5) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_46 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(n11), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI22_X1 U4 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U8 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U10 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U11 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U16 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U17 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U18 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U19 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U20 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U21 ( .A(Ci), .ZN(n46) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_47 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n7) );
  INV_X1 U2 ( .A(n12), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI22_X1 U4 ( .A1(n9), .A2(n1), .B1(Ci), .B2(n8), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n10), .A2(n7), .B1(n5), .B2(n4), .ZN(n9) );
  AOI22_X1 U6 ( .A1(n7), .A2(n30), .B1(n6), .B2(n5), .ZN(n8) );
  NAND2_X1 U7 ( .A1(n3), .A2(n13), .ZN(n5) );
  OAI22_X1 U8 ( .A1(n36), .A2(n1), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(n37), .A2(n34), .B1(n33), .B2(n12), .ZN(n36) );
  AOI22_X1 U10 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U11 ( .A1(n11), .A2(n39), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n1), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U16 ( .A(Ci), .B(n2), .ZN(S[0]) );
  NAND2_X1 U17 ( .A1(n4), .A2(n30), .ZN(n2) );
  OAI21_X1 U18 ( .B1(n31), .B2(n30), .A(n13), .ZN(n32) );
  OAI21_X1 U19 ( .B1(n10), .B2(n31), .A(n13), .ZN(n12) );
  OAI21_X1 U20 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U21 ( .A(n10), .ZN(n4) );
  INV_X1 U22 ( .A(n30), .ZN(n6) );
  INV_X1 U23 ( .A(n40), .ZN(n11) );
  INV_X1 U24 ( .A(n31), .ZN(n3) );
  NOR2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U29 ( .A1(B[1]), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  INV_X1 U31 ( .A(Ci), .ZN(n1) );
endmodule


module carry_sel_bk_NB4_49 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
endmodule


module carry_sel_bk_NB4_50 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U11 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U12 ( .A(n30), .ZN(n5) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
endmodule


module carry_sel_bk_NB4_51 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n40), .ZN(n10) );
  INV_X1 U24 ( .A(n30), .ZN(n5) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NAND2_X1 U27 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_55 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(n11), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI21_X1 U4 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U5 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U6 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U7 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U8 ( .A(n31), .ZN(n2) );
  INV_X1 U9 ( .A(n9), .ZN(n3) );
  INV_X1 U10 ( .A(n40), .ZN(n10) );
  OAI22_X1 U11 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U12 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U13 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U14 ( .A(n30), .ZN(n5) );
  OAI22_X1 U15 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U16 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U17 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U18 ( .A1(n10), .A2(n39), .ZN(n33) );
  XNOR2_X1 U19 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U20 ( .A1(n3), .A2(n30), .ZN(n1) );
  NOR2_X1 U21 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U22 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  OAI22_X1 U23 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U24 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U25 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U26 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  INV_X1 U27 ( .A(Ci), .ZN(n46) );
  NAND2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U29 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NOR2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_58 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NOR2_X1 U28 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_59 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  AOI22_X1 U7 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  INV_X1 U8 ( .A(n30), .ZN(n5) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  NAND2_X1 U22 ( .A1(n2), .A2(n12), .ZN(n4) );
  INV_X1 U23 ( .A(n31), .ZN(n2) );
  INV_X1 U24 ( .A(n9), .ZN(n3) );
  INV_X1 U25 ( .A(n40), .ZN(n10) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NAND2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U30 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
endmodule


module carry_sel_bk_NB4_61 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U9 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U11 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module carry_sel_bk_NB4_62 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(Ci), .ZN(n46) );
  INV_X1 U3 ( .A(n11), .ZN(n37) );
  INV_X1 U4 ( .A(n32), .ZN(n41) );
  OAI22_X1 U5 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U6 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U7 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U8 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U9 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U13 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U14 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U15 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U16 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U17 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U18 ( .A1(n3), .A2(n30), .ZN(n1) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n30), .ZN(n5) );
  INV_X1 U24 ( .A(n40), .ZN(n10) );
  INV_X1 U25 ( .A(n31), .ZN(n2) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
endmodule


module carry_sel_bk_NB4_63 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n42) );
  XOR2_X1 U33 ( .A(A[2]), .B(B[2]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[1]), .B(B[1]), .Z(n6) );
  INV_X1 U2 ( .A(n11), .ZN(n37) );
  INV_X1 U3 ( .A(n32), .ZN(n41) );
  OAI22_X1 U4 ( .A1(n8), .A2(n46), .B1(Ci), .B2(n7), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(n9), .A2(n6), .B1(n4), .B2(n3), .ZN(n8) );
  AOI22_X1 U6 ( .A1(n6), .A2(n30), .B1(n5), .B2(n4), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n2), .A2(n12), .ZN(n4) );
  OAI22_X1 U8 ( .A1(n36), .A2(n46), .B1(Ci), .B2(n35), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(n37), .A2(n34), .B1(n33), .B2(n11), .ZN(n36) );
  AOI22_X1 U10 ( .A1(n41), .A2(n34), .B1(n33), .B2(n32), .ZN(n35) );
  NAND2_X1 U11 ( .A1(n10), .A2(n39), .ZN(n33) );
  OAI22_X1 U12 ( .A1(n46), .A2(n45), .B1(Ci), .B2(n44), .ZN(S[3]) );
  XNOR2_X1 U13 ( .A(n43), .B(n42), .ZN(n44) );
  XNOR2_X1 U14 ( .A(n38), .B(n42), .ZN(n45) );
  OAI21_X1 U15 ( .B1(n41), .B2(n40), .A(n39), .ZN(n43) );
  XNOR2_X1 U16 ( .A(Ci), .B(n1), .ZN(S[0]) );
  NAND2_X1 U17 ( .A1(n3), .A2(n30), .ZN(n1) );
  INV_X1 U18 ( .A(Ci), .ZN(n46) );
  OAI21_X1 U19 ( .B1(n31), .B2(n30), .A(n12), .ZN(n32) );
  OAI21_X1 U20 ( .B1(n9), .B2(n31), .A(n12), .ZN(n11) );
  OAI21_X1 U21 ( .B1(n37), .B2(n40), .A(n39), .ZN(n38) );
  INV_X1 U22 ( .A(n9), .ZN(n3) );
  INV_X1 U23 ( .A(n40), .ZN(n10) );
  INV_X1 U24 ( .A(n31), .ZN(n2) );
  INV_X1 U25 ( .A(n30), .ZN(n5) );
  NOR2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n31) );
  NOR2_X1 U28 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(A[0]), .ZN(n30) );
  NAND2_X1 U30 ( .A1(B[1]), .A2(A[1]), .ZN(n12) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
endmodule


module sum_gen_Nrca4_NB32_0 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_7 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  carry_sel_bk_NB4_6 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  carry_sel_bk_NB4_5 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  carry_sel_bk_NB4_4 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_3 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_2 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_1 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_0 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_0 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_31 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_30 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_29 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_28 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_27 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_26 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_25 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_24 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_23 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_22 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_21 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_20 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_19 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_18 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_17 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_16 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_15 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_14 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_13 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_12 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_11 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_10 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_9 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_8 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_7 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_6 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_5 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_4 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_3 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_2 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_1 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_0 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_26 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_8 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_25 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_24 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_23 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_22 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_21 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_20 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_19 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_18 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_17 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_16 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_15 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_14 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_13 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_12 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_7 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_11 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_10 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_9 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_8 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_7 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_6 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_5 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_6 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_4 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_3 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_2 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_5 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_4 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_1 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_0 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_3 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_2 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_1 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_0 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module sum_gen_Nrca4_NB32_1 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_15 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_14 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_13 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_12 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_11 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_10 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_9 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_8 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_1 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_63 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_62 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_61 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_60 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_59 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_58 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_57 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_56 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_55 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_54 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_53 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_52 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_51 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_50 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_49 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_48 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_47 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_46 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_45 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_44 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_43 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_42 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_41 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_40 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_39 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_38 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_37 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_36 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_35 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_34 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_33 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_32 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_53 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_17 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_52 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_51 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_50 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_49 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_48 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_47 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_46 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_45 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_44 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_43 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_42 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_41 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_40 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_39 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_16 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_38 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_37 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_36 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_35 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_34 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_33 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_32 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_15 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_31 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_30 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_29 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_14 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_13 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_28 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_27 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_12 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_11 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_10 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_9 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module sum_gen_Nrca4_NB32_2 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_23 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_22 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_21 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_20 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_19 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_18 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_17 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_16 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_3 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_31 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_30 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_29 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_28 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_27 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_26 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_25 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_24 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_3 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_127 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_126 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_125 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_124 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_123 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_122 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_121 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_120 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_119 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_118 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_117 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_116 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_115 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_114 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_113 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_112 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_111 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_110 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_109 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_108 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_107 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_106 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_105 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_104 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_103 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_102 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_101 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_100 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_99 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_98 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_97 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_96 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_107 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_35 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_106 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_105 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_104 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_103 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_102 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_101 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_100 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_99 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_98 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_97 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_96 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_95 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_94 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_93 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_34 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_92 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_91 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_90 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_89 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_88 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_87 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_86 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_33 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_85 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_84 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_83 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_32 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_31 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_82 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_81 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_30 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_29 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_28 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_27 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module sum_gen_Nrca4_NB32_4 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_39 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_38 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_37 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_36 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_35 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_34 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_33 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_32 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_5 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_47 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_46 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_45 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_44 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_43 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_42 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_41 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_40 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_6 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_55 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_54 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_53 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_52 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_51 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_50 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_49 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_48 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_7 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_63 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_62 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_61 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_60 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_59 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_58 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_57 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_56 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_7 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1;

  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(\matrixGen[0][0] ) );
  pg_net_255 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_254 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_253 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_252 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_251 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_250 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_249 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_248 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_247 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_246 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_245 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_244 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_243 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_242 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_241 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_240 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_239 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_238 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_237 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_236 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_235 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_234 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_233 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_232 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_231 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_230 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_229 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_228 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_227 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_226 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_225 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_224 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_215 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_71 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_214 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_213 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_212 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_211 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_210 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_209 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_208 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_207 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_206 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_205 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_204 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_203 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_202 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_201 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_70 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_200 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_199 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_198 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_197 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_196 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_195 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_194 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_69 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_193 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_192 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_191 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_68 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_67 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_190 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_189 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_66 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_65 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_64 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_63 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
endmodule


module carry_sel_bk_NB4_64 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32;

  XNOR2_X1 U3 ( .A(n24), .B(n3), .ZN(n28) );
  XNOR2_X1 U4 ( .A(n3), .B(n26), .ZN(n27) );
  OAI21_X1 U5 ( .B1(n20), .B2(n19), .A(n18), .ZN(n25) );
  OAI21_X1 U6 ( .B1(n20), .B2(n16), .A(n18), .ZN(n23) );
  NAND2_X1 U7 ( .A1(n8), .A2(n9), .ZN(n17) );
  NAND2_X1 U9 ( .A1(A[0]), .A2(B[0]), .ZN(n16) );
  NAND2_X1 U10 ( .A1(A[1]), .A2(B[1]), .ZN(n18) );
  NOR2_X1 U11 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  AND2_X1 U12 ( .A1(A[2]), .A2(B[2]), .ZN(n2) );
  XOR2_X1 U13 ( .A(A[3]), .B(B[3]), .Z(n3) );
  XOR2_X1 U14 ( .A(B[2]), .B(A[2]), .Z(n22) );
  OR2_X1 U15 ( .A1(B[2]), .A2(A[2]), .ZN(n4) );
  INV_X1 U16 ( .A(A[0]), .ZN(n8) );
  INV_X1 U17 ( .A(B[0]), .ZN(n9) );
  NAND2_X1 U18 ( .A1(n16), .A2(n17), .ZN(n5) );
  NAND2_X1 U20 ( .A1(Ci), .A2(n17), .ZN(n6) );
  NAND2_X1 U21 ( .A1(n16), .A2(n6), .ZN(n15) );
  NAND2_X1 U22 ( .A1(Ci), .A2(B[0]), .ZN(n7) );
  NAND2_X1 U23 ( .A1(n7), .A2(n8), .ZN(n12) );
  INV_X1 U24 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U25 ( .A1(n10), .A2(n9), .ZN(n11) );
  NAND2_X1 U26 ( .A1(n12), .A2(n11), .ZN(n14) );
  INV_X1 U27 ( .A(A[1]), .ZN(n13) );
  INV_X1 U28 ( .A(n17), .ZN(n19) );
  OAI21_X1 U29 ( .B1(n23), .B2(Ci), .A(n25), .ZN(n21) );
  XNOR2_X1 U30 ( .A(n21), .B(n22), .ZN(S[2]) );
  AOI21_X1 U31 ( .B1(n23), .B2(n4), .A(n2), .ZN(n24) );
  AOI21_X1 U32 ( .B1(n25), .B2(n4), .A(n2), .ZN(n26) );
  MUX2_X1 U33 ( .A(n28), .B(n27), .S(n32), .Z(S[3]) );
  NAND2_X1 U2 ( .A1(n14), .A2(n29), .ZN(n30) );
  NAND2_X2 U8 ( .A1(n15), .A2(n1), .ZN(n31) );
  NAND2_X1 U19 ( .A1(n30), .A2(n31), .ZN(S[1]) );
  INV_X1 U34 ( .A(n1), .ZN(n29) );
  XOR2_X2 U35 ( .A(B[1]), .B(n13), .Z(n1) );
  XNOR2_X2 U36 ( .A(n32), .B(n5), .ZN(S[0]) );
  BUF_X1 U37 ( .A(Ci), .Z(n32) );
endmodule


module carry_sel_bk_NB4_65 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32;

  XOR2_X1 U2 ( .A(B[1]), .B(n17), .Z(n8) );
  INV_X1 U3 ( .A(n8), .ZN(n2) );
  XOR2_X1 U4 ( .A(A[3]), .B(B[3]), .Z(n1) );
  NAND2_X1 U5 ( .A1(n18), .A2(n2), .ZN(n3) );
  NAND2_X1 U6 ( .A1(n19), .A2(n8), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n3), .A2(n4), .ZN(S[1]) );
  XNOR2_X1 U9 ( .A(n28), .B(n1), .ZN(n32) );
  XNOR2_X1 U10 ( .A(n1), .B(n30), .ZN(n31) );
  OAI21_X1 U11 ( .B1(n24), .B2(n23), .A(n22), .ZN(n29) );
  OAI21_X1 U12 ( .B1(n24), .B2(n20), .A(n22), .ZN(n27) );
  NAND2_X1 U13 ( .A1(n12), .A2(n13), .ZN(n21) );
  XOR2_X1 U14 ( .A(B[2]), .B(A[2]), .Z(n26) );
  NAND2_X1 U15 ( .A1(A[1]), .A2(B[1]), .ZN(n22) );
  NAND2_X1 U16 ( .A1(A[0]), .A2(B[0]), .ZN(n20) );
  NOR2_X1 U17 ( .A1(B[1]), .A2(A[1]), .ZN(n24) );
  AND2_X1 U18 ( .A1(A[2]), .A2(B[2]), .ZN(n6) );
  OR2_X1 U19 ( .A1(B[2]), .A2(A[2]), .ZN(n7) );
  INV_X1 U20 ( .A(A[0]), .ZN(n12) );
  INV_X1 U21 ( .A(B[0]), .ZN(n13) );
  NAND2_X1 U22 ( .A1(n20), .A2(n21), .ZN(n9) );
  XNOR2_X1 U23 ( .A(Ci), .B(n9), .ZN(S[0]) );
  NAND2_X1 U24 ( .A1(Ci), .A2(n21), .ZN(n10) );
  NAND2_X1 U25 ( .A1(n20), .A2(n10), .ZN(n19) );
  NAND2_X1 U26 ( .A1(Ci), .A2(B[0]), .ZN(n11) );
  NAND2_X1 U27 ( .A1(n11), .A2(n12), .ZN(n16) );
  INV_X1 U28 ( .A(Ci), .ZN(n14) );
  NAND2_X1 U29 ( .A1(n14), .A2(n13), .ZN(n15) );
  NAND2_X1 U30 ( .A1(n16), .A2(n15), .ZN(n18) );
  INV_X1 U31 ( .A(A[1]), .ZN(n17) );
  INV_X1 U32 ( .A(n21), .ZN(n23) );
  OAI21_X1 U33 ( .B1(Ci), .B2(n27), .A(n29), .ZN(n25) );
  XNOR2_X1 U34 ( .A(n25), .B(n26), .ZN(S[2]) );
  AOI21_X1 U35 ( .B1(n27), .B2(n7), .A(n6), .ZN(n28) );
  AOI21_X1 U36 ( .B1(n29), .B2(n7), .A(n6), .ZN(n30) );
  MUX2_X1 U37 ( .A(n32), .B(n31), .S(Ci), .Z(S[3]) );
endmodule


module carry_sel_bk_NB4_66 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45;

  XOR2_X1 U2 ( .A(A[3]), .B(B[3]), .Z(n1) );
  XNOR2_X1 U5 ( .A(n25), .B(n1), .ZN(n29) );
  XNOR2_X1 U6 ( .A(n1), .B(n27), .ZN(n28) );
  OAI21_X1 U7 ( .B1(n21), .B2(n20), .A(n19), .ZN(n26) );
  XOR2_X1 U13 ( .A(B[2]), .B(A[2]), .Z(n23) );
  AND2_X1 U14 ( .A1(A[2]), .A2(B[2]), .ZN(n3) );
  OR2_X1 U15 ( .A1(B[2]), .A2(A[2]), .ZN(n4) );
  XNOR2_X1 U19 ( .A(n2), .B(n5), .ZN(S[0]) );
  OAI21_X1 U30 ( .B1(n24), .B2(Ci), .A(n26), .ZN(n22) );
  XNOR2_X1 U31 ( .A(n22), .B(n23), .ZN(S[2]) );
  AOI21_X1 U32 ( .B1(n24), .B2(n4), .A(n3), .ZN(n25) );
  AOI21_X1 U33 ( .B1(n26), .B2(n4), .A(n3), .ZN(n27) );
  MUX2_X1 U34 ( .A(n29), .B(n28), .S(Ci), .Z(S[3]) );
  NAND2_X2 syn91 ( .A1(n44), .A2(n43), .ZN(n33) );
  INV_X2 syn90 ( .A(n19), .ZN(n38) );
  INV_X2 syn87 ( .A(n32), .ZN(n44) );
  INV_X2 syn63 ( .A(n43), .ZN(n21) );
  NAND2_X2 syn62 ( .A1(n36), .A2(n37), .ZN(n43) );
  INV_X2 syn58 ( .A(n31), .ZN(n20) );
  NAND2_X2 syn57 ( .A1(n34), .A2(n35), .ZN(n31) );
  INV_X2 syn20 ( .A(A[1]), .ZN(n36) );
  INV_X2 syn14 ( .A(A[0]), .ZN(n35) );
  INV_X2 syn13 ( .A(B[0]), .ZN(n34) );
  NAND2_X2 syn10 ( .A1(A[0]), .A2(B[0]), .ZN(n32) );
  NAND2_X2 net432328 ( .A1(n19), .A2(n33), .ZN(n24) );
  NAND2_X2 net432330 ( .A1(n31), .A2(n32), .ZN(n5) );
  MUX2_X2 U3 ( .A(n41), .B(n40), .S(n30), .Z(S[1]) );
  OR2_X1 U4 ( .A1(n38), .A2(n21), .ZN(n30) );
  NAND2_X1 U8 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  INV_X1 U9 ( .A(B[1]), .ZN(n37) );
  INV_X1 U10 ( .A(Ci), .ZN(n39) );
  INV_X1 U11 ( .A(n39), .ZN(n2) );
  NAND2_X1 U12 ( .A1(n32), .A2(n45), .ZN(n42) );
  OAI21_X1 U16 ( .B1(n20), .B2(n39), .A(n32), .ZN(n40) );
  INV_X1 U17 ( .A(Ci), .ZN(n45) );
  NAND2_X1 U18 ( .A1(n42), .A2(n31), .ZN(n41) );
endmodule


module carry_sel_bk_NB4_67 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  XOR2_X1 U2 ( .A(A[3]), .B(B[3]), .Z(n1) );
  XNOR2_X1 U3 ( .A(n24), .B(n1), .ZN(n28) );
  XNOR2_X1 U4 ( .A(n1), .B(n26), .ZN(n27) );
  OAI21_X1 U5 ( .B1(n20), .B2(n19), .A(n18), .ZN(n25) );
  OAI21_X1 U6 ( .B1(n20), .B2(n16), .A(n18), .ZN(n23) );
  NAND2_X1 U7 ( .A1(n8), .A2(n9), .ZN(n17) );
  MUX2_X1 U8 ( .A(n14), .B(n15), .S(n2), .Z(S[1]) );
  XOR2_X1 U9 ( .A(B[1]), .B(n13), .Z(n2) );
  XOR2_X1 U10 ( .A(B[2]), .B(A[2]), .Z(n22) );
  NAND2_X1 U11 ( .A1(A[0]), .A2(B[0]), .ZN(n16) );
  AND2_X1 U12 ( .A1(A[2]), .A2(B[2]), .ZN(n3) );
  OR2_X1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n4) );
  NAND2_X1 U14 ( .A1(A[1]), .A2(B[1]), .ZN(n18) );
  NOR2_X1 U15 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  INV_X1 U16 ( .A(A[0]), .ZN(n8) );
  INV_X1 U17 ( .A(B[0]), .ZN(n9) );
  NAND2_X1 U18 ( .A1(n16), .A2(n17), .ZN(n5) );
  XNOR2_X1 U19 ( .A(Ci), .B(n5), .ZN(S[0]) );
  NAND2_X1 U20 ( .A1(Ci), .A2(n17), .ZN(n6) );
  NAND2_X1 U21 ( .A1(n16), .A2(n6), .ZN(n15) );
  NAND2_X1 U22 ( .A1(Ci), .A2(B[0]), .ZN(n7) );
  NAND2_X1 U23 ( .A1(n8), .A2(n7), .ZN(n12) );
  INV_X1 U24 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U25 ( .A1(n10), .A2(n9), .ZN(n11) );
  NAND2_X1 U26 ( .A1(n12), .A2(n11), .ZN(n14) );
  INV_X1 U27 ( .A(A[1]), .ZN(n13) );
  INV_X1 U28 ( .A(n17), .ZN(n19) );
  OAI21_X1 U29 ( .B1(n23), .B2(Ci), .A(n25), .ZN(n21) );
  XNOR2_X1 U30 ( .A(n22), .B(n21), .ZN(S[2]) );
  AOI21_X1 U31 ( .B1(n23), .B2(n4), .A(n3), .ZN(n24) );
  AOI21_X1 U32 ( .B1(n25), .B2(n4), .A(n3), .ZN(n26) );
  MUX2_X1 U33 ( .A(n28), .B(n27), .S(Ci), .Z(S[3]) );
endmodule


module carry_sel_bk_NB4_68 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  XOR2_X1 U2 ( .A(A[3]), .B(B[3]), .Z(n1) );
  OAI21_X1 U3 ( .B1(n24), .B2(n23), .A(n22), .ZN(n28) );
  MUX2_X1 U4 ( .A(n18), .B(n19), .S(n2), .Z(S[1]) );
  XOR2_X1 U5 ( .A(B[1]), .B(n8), .Z(n2) );
  XNOR2_X1 U6 ( .A(n27), .B(n1), .ZN(n31) );
  XNOR2_X1 U7 ( .A(n1), .B(n29), .ZN(n30) );
  OAI21_X1 U8 ( .B1(n24), .B2(n20), .A(n22), .ZN(n26) );
  NAND2_X1 U9 ( .A1(n6), .A2(n14), .ZN(n21) );
  XOR2_X1 U10 ( .A(n3), .B(n25), .Z(S[2]) );
  XOR2_X1 U11 ( .A(B[2]), .B(n10), .Z(n3) );
  OR2_X1 U12 ( .A1(B[2]), .A2(n9), .ZN(n4) );
  AND2_X1 U13 ( .A1(n9), .A2(B[2]), .ZN(n5) );
  NAND2_X1 U14 ( .A1(n7), .A2(B[1]), .ZN(n22) );
  NOR2_X1 U15 ( .A1(B[1]), .A2(n7), .ZN(n24) );
  NAND2_X1 U16 ( .A1(A[0]), .A2(B[0]), .ZN(n20) );
  INV_X1 U17 ( .A(A[0]), .ZN(n6) );
  INV_X1 U18 ( .A(n8), .ZN(n7) );
  INV_X1 U19 ( .A(A[1]), .ZN(n8) );
  INV_X1 U20 ( .A(n10), .ZN(n9) );
  INV_X1 U21 ( .A(A[2]), .ZN(n10) );
  INV_X1 U22 ( .A(B[0]), .ZN(n14) );
  NAND2_X1 U23 ( .A1(n20), .A2(n21), .ZN(n11) );
  XNOR2_X1 U24 ( .A(Ci), .B(n11), .ZN(S[0]) );
  NAND2_X1 U25 ( .A1(Ci), .A2(n21), .ZN(n12) );
  NAND2_X1 U26 ( .A1(n20), .A2(n12), .ZN(n19) );
  NAND2_X1 U27 ( .A1(Ci), .A2(B[0]), .ZN(n13) );
  NAND2_X1 U28 ( .A1(n6), .A2(n13), .ZN(n17) );
  INV_X1 U29 ( .A(Ci), .ZN(n15) );
  NAND2_X1 U30 ( .A1(n15), .A2(n14), .ZN(n16) );
  NAND2_X1 U31 ( .A1(n17), .A2(n16), .ZN(n18) );
  INV_X1 U32 ( .A(n21), .ZN(n23) );
  OAI21_X1 U33 ( .B1(n26), .B2(Ci), .A(n28), .ZN(n25) );
  AOI21_X1 U34 ( .B1(n26), .B2(n4), .A(n5), .ZN(n27) );
  AOI21_X1 U35 ( .B1(n28), .B2(n4), .A(n5), .ZN(n29) );
  MUX2_X1 U36 ( .A(n31), .B(n30), .S(Ci), .Z(S[3]) );
endmodule


module carry_sel_bk_NB4_69 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  XOR2_X1 U2 ( .A(A[3]), .B(B[3]), .Z(n1) );
  OAI21_X1 U3 ( .B1(n23), .B2(n22), .A(n21), .ZN(n28) );
  OAI21_X1 U4 ( .B1(n23), .B2(n19), .A(n21), .ZN(n26) );
  XNOR2_X1 U5 ( .A(n27), .B(n1), .ZN(n31) );
  XNOR2_X1 U6 ( .A(n1), .B(n29), .ZN(n30) );
  NAND2_X1 U7 ( .A1(n5), .A2(n13), .ZN(n20) );
  OR2_X1 U8 ( .A1(B[2]), .A2(n8), .ZN(n2) );
  AND2_X1 U9 ( .A1(n8), .A2(B[2]), .ZN(n3) );
  MUX2_X1 U10 ( .A(n17), .B(n18), .S(n4), .Z(S[1]) );
  XOR2_X1 U11 ( .A(B[1]), .B(n7), .Z(n4) );
  NAND2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n19) );
  NAND2_X1 U13 ( .A1(n6), .A2(B[1]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(n6), .ZN(n23) );
  INV_X1 U15 ( .A(A[0]), .ZN(n5) );
  INV_X1 U16 ( .A(n7), .ZN(n6) );
  INV_X1 U17 ( .A(A[1]), .ZN(n7) );
  INV_X1 U18 ( .A(n9), .ZN(n8) );
  INV_X1 U19 ( .A(A[2]), .ZN(n9) );
  INV_X1 U20 ( .A(B[0]), .ZN(n13) );
  NAND2_X1 U21 ( .A1(n19), .A2(n20), .ZN(n10) );
  XNOR2_X1 U22 ( .A(Ci), .B(n10), .ZN(S[0]) );
  NAND2_X1 U23 ( .A1(Ci), .A2(n20), .ZN(n11) );
  NAND2_X1 U24 ( .A1(n19), .A2(n11), .ZN(n18) );
  NAND2_X1 U25 ( .A1(Ci), .A2(B[0]), .ZN(n12) );
  NAND2_X1 U26 ( .A1(n5), .A2(n12), .ZN(n16) );
  INV_X1 U27 ( .A(Ci), .ZN(n14) );
  NAND2_X1 U28 ( .A1(n14), .A2(n13), .ZN(n15) );
  NAND2_X1 U29 ( .A1(n16), .A2(n15), .ZN(n17) );
  XNOR2_X1 U30 ( .A(B[2]), .B(n9), .ZN(n25) );
  INV_X1 U31 ( .A(n20), .ZN(n22) );
  OAI21_X1 U32 ( .B1(n26), .B2(Ci), .A(n28), .ZN(n24) );
  XNOR2_X1 U33 ( .A(n25), .B(n24), .ZN(S[2]) );
  AOI21_X1 U34 ( .B1(n26), .B2(n2), .A(n3), .ZN(n27) );
  AOI21_X1 U35 ( .B1(n28), .B2(n2), .A(n3), .ZN(n29) );
  MUX2_X1 U36 ( .A(n31), .B(n30), .S(Ci), .Z(S[3]) );
endmodule


module carry_sel_bk_NB4_70 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  XOR2_X1 U2 ( .A(A[3]), .B(B[3]), .Z(n1) );
  XNOR2_X1 U3 ( .A(n27), .B(n1), .ZN(n31) );
  XNOR2_X1 U4 ( .A(n1), .B(n29), .ZN(n30) );
  OAI21_X1 U5 ( .B1(n23), .B2(n19), .A(n21), .ZN(n26) );
  OAI21_X1 U6 ( .B1(n23), .B2(n22), .A(n21), .ZN(n28) );
  NAND2_X1 U7 ( .A1(n5), .A2(n13), .ZN(n20) );
  OR2_X1 U8 ( .A1(B[2]), .A2(n8), .ZN(n2) );
  AND2_X1 U9 ( .A1(n8), .A2(B[2]), .ZN(n3) );
  MUX2_X1 U10 ( .A(n17), .B(n18), .S(n4), .Z(S[1]) );
  XOR2_X1 U11 ( .A(B[1]), .B(n7), .Z(n4) );
  NAND2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n19) );
  NAND2_X1 U13 ( .A1(n6), .A2(B[1]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(n6), .ZN(n23) );
  INV_X1 U15 ( .A(A[0]), .ZN(n5) );
  INV_X1 U16 ( .A(n7), .ZN(n6) );
  INV_X1 U17 ( .A(A[1]), .ZN(n7) );
  INV_X1 U18 ( .A(n9), .ZN(n8) );
  INV_X1 U19 ( .A(A[2]), .ZN(n9) );
  INV_X1 U20 ( .A(B[0]), .ZN(n13) );
  NAND2_X1 U21 ( .A1(n19), .A2(n20), .ZN(n10) );
  XNOR2_X1 U22 ( .A(Ci), .B(n10), .ZN(S[0]) );
  NAND2_X1 U23 ( .A1(Ci), .A2(n20), .ZN(n11) );
  NAND2_X1 U24 ( .A1(n19), .A2(n11), .ZN(n18) );
  NAND2_X1 U25 ( .A1(Ci), .A2(B[0]), .ZN(n12) );
  NAND2_X1 U26 ( .A1(n5), .A2(n12), .ZN(n16) );
  INV_X1 U27 ( .A(Ci), .ZN(n14) );
  NAND2_X1 U28 ( .A1(n14), .A2(n13), .ZN(n15) );
  NAND2_X1 U29 ( .A1(n16), .A2(n15), .ZN(n17) );
  XNOR2_X1 U30 ( .A(B[2]), .B(n9), .ZN(n25) );
  INV_X1 U31 ( .A(n20), .ZN(n22) );
  OAI21_X1 U32 ( .B1(n26), .B2(Ci), .A(n28), .ZN(n24) );
  XNOR2_X1 U33 ( .A(n25), .B(n24), .ZN(S[2]) );
  AOI21_X1 U34 ( .B1(n26), .B2(n2), .A(n3), .ZN(n27) );
  AOI21_X1 U35 ( .B1(n28), .B2(n2), .A(n3), .ZN(n29) );
  MUX2_X1 U36 ( .A(n31), .B(n30), .S(Ci), .Z(S[3]) );
endmodule


module carry_sel_bk_NB4_71 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  XOR2_X1 U2 ( .A(A[3]), .B(B[3]), .Z(n1) );
  OAI21_X1 U3 ( .B1(n22), .B2(n21), .A(n20), .ZN(n27) );
  OR2_X1 U4 ( .A1(B[2]), .A2(A[2]), .ZN(n2) );
  AND2_X1 U5 ( .A1(A[2]), .A2(B[2]), .ZN(n3) );
  XOR2_X1 U6 ( .A(n10), .B(n4), .Z(S[0]) );
  AND2_X1 U7 ( .A1(n19), .A2(n12), .ZN(n4) );
  XNOR2_X1 U8 ( .A(n26), .B(n1), .ZN(n30) );
  XNOR2_X1 U9 ( .A(n1), .B(n28), .ZN(n29) );
  OAI21_X1 U10 ( .B1(n22), .B2(n19), .A(n20), .ZN(n25) );
  NAND2_X1 U11 ( .A1(n6), .A2(n14), .ZN(n12) );
  MUX2_X1 U12 ( .A(n17), .B(n18), .S(n5), .Z(S[1]) );
  XOR2_X1 U13 ( .A(B[1]), .B(n8), .Z(n5) );
  NAND2_X1 U14 ( .A1(A[0]), .A2(B[0]), .ZN(n19) );
  NAND2_X1 U15 ( .A1(n7), .A2(B[1]), .ZN(n20) );
  NOR2_X1 U16 ( .A1(B[1]), .A2(n7), .ZN(n22) );
  INV_X1 U17 ( .A(A[0]), .ZN(n6) );
  INV_X1 U18 ( .A(n8), .ZN(n7) );
  INV_X1 U19 ( .A(A[1]), .ZN(n8) );
  INV_X1 U20 ( .A(A[2]), .ZN(n9) );
  INV_X1 U21 ( .A(n11), .ZN(n10) );
  INV_X1 U22 ( .A(Ci), .ZN(n11) );
  INV_X1 U23 ( .A(B[0]), .ZN(n14) );
  INV_X1 U24 ( .A(n12), .ZN(n21) );
  OAI21_X1 U25 ( .B1(n21), .B2(n11), .A(n19), .ZN(n18) );
  NAND2_X1 U26 ( .A1(n10), .A2(B[0]), .ZN(n13) );
  NAND2_X1 U27 ( .A1(n6), .A2(n13), .ZN(n16) );
  NAND2_X1 U28 ( .A1(n11), .A2(n14), .ZN(n15) );
  NAND2_X1 U29 ( .A1(n16), .A2(n15), .ZN(n17) );
  XNOR2_X1 U30 ( .A(B[2]), .B(n9), .ZN(n24) );
  OAI21_X1 U31 ( .B1(n25), .B2(n10), .A(n27), .ZN(n23) );
  XNOR2_X1 U32 ( .A(n24), .B(n23), .ZN(S[2]) );
  AOI21_X1 U33 ( .B1(n25), .B2(n2), .A(n3), .ZN(n26) );
  AOI21_X1 U34 ( .B1(n27), .B2(n2), .A(n3), .ZN(n28) );
  MUX2_X1 U35 ( .A(n30), .B(n29), .S(n10), .Z(S[3]) );
endmodule


module G_72 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2, n1;

  INV_X1 U2 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U1 ( .A1(Gk_1j), .A2(Pik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n1), .A2(n2), .ZN(Gij) );
endmodule


module G_73 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1, n2;

  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(Gij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n1) );
  INV_X1 U3 ( .A(Gik), .ZN(n2) );
endmodule


module G_74 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1, n2;

  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n1) );
  INV_X1 U3 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Gij) );
endmodule


module G_75 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n1) );
endmodule


module blockPG_217 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module G_76 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(Gk_1j), .A2(Pik), .ZN(n1) );
  INV_X1 U2 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(Gij) );
endmodule


module G_77 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2, n1;

  INV_X1 U3 ( .A(Gik), .ZN(n2) );
  NAND2_X2 U1 ( .A1(n2), .A2(n1), .ZN(Gij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n1) );
endmodule


module blockPG_218 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module blockPG_220 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module G_79 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2, n1;

  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n1) );
  INV_X1 U3 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_229 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_232 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  OR2_X1 U2 ( .A1(Gik), .A2(n2), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
endmodule


module blockPG_233 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  NAND2_X1 U1 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_237 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_238 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module blockPG_239 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Gk_1j), .A2(Pik), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module blockPG_241 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module G_80 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(Gk_1j), .A2(Pik), .ZN(n1) );
  INV_X1 U2 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n1), .A2(n2), .ZN(Gij) );
endmodule


module blockPG_242 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2, n3;

  AND2_X1 U1 ( .A1(Pik), .A2(Pk_1j), .ZN(Pij) );
  NAND2_X1 U2 ( .A1(Pik), .A2(Gk_1j), .ZN(n2) );
  INV_X1 U3 ( .A(Gik), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(Gij) );
endmodule


module pg_net_259 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_280 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module pg_net_282 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_283 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p) );
endmodule


module pg_net_284 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module pg_net_286 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module pg_net_287 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module p4addgen_NB32_CW4_0 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_0 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_0 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_1 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_1 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_1 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_2 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_2 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_2 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_3 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_3 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_3 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_4 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_4 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_4 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_5 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_5 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_5 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_6 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_6 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_6 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_7 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_7 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_7 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module MUX_SHIFT_NB16_N_sh14_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   \B[30] , \B[0] , n63, n2, n3, n4, n5, n6, n1, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n62;
  assign B[31] = \B[30] ;
  assign B[30] = \B[30] ;
  assign AS = \B[0] ;
  assign B[13] = \B[0] ;
  assign B[12] = \B[0] ;
  assign B[11] = \B[0] ;
  assign B[10] = \B[0] ;
  assign B[9] = \B[0] ;
  assign B[8] = \B[0] ;
  assign B[7] = \B[0] ;
  assign B[6] = \B[0] ;
  assign B[5] = \B[0] ;
  assign B[4] = \B[0] ;
  assign B[3] = \B[0] ;
  assign B[2] = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  CLKBUF_X3 U3 ( .A(n63), .Z(\B[0] ) );
  XOR2_X2 U4 ( .A(n12), .B(sel[2]), .Z(n11) );
  XNOR2_X1 U5 ( .A(n12), .B(sel[0]), .ZN(n7) );
  XNOR2_X1 U6 ( .A(n12), .B(sel[0]), .ZN(n1) );
  XNOR2_X1 U7 ( .A(n12), .B(sel[0]), .ZN(n8) );
  INV_X1 U8 ( .A(n2), .ZN(B[14]) );
  AOI22_X1 U9 ( .A1(n3), .A2(\B[0] ), .B1(n4), .B2(n5), .ZN(n2) );
  INV_X1 U10 ( .A(n3), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  NOR2_X1 U12 ( .A1(n20), .A2(n11), .ZN(n45) );
  NOR2_X1 U13 ( .A1(n18), .A2(n11), .ZN(n44) );
  NOR2_X1 U14 ( .A1(n28), .A2(n11), .ZN(n49) );
  NOR2_X1 U15 ( .A1(n26), .A2(n11), .ZN(n48) );
  NOR2_X1 U16 ( .A1(n36), .A2(n11), .ZN(n53) );
  NOR2_X1 U17 ( .A1(n34), .A2(n11), .ZN(n52) );
  NOR2_X1 U18 ( .A1(n41), .A2(n11), .ZN(n56) );
  NOR2_X1 U19 ( .A1(n16), .A2(n11), .ZN(n43) );
  NOR2_X1 U20 ( .A1(n24), .A2(n11), .ZN(n47) );
  NOR2_X1 U21 ( .A1(n32), .A2(n11), .ZN(n51) );
  NOR2_X1 U22 ( .A1(n40), .A2(n11), .ZN(n55) );
  INV_X1 U23 ( .A(n59), .ZN(\B[30] ) );
  NAND2_X1 U24 ( .A1(n9), .A2(n57), .ZN(n58) );
  NOR2_X1 U25 ( .A1(n11), .A2(n13), .ZN(n42) );
  NOR2_X1 U27 ( .A1(n38), .A2(n11), .ZN(n54) );
  NOR2_X1 U28 ( .A1(n30), .A2(n11), .ZN(n50) );
  NOR2_X1 U29 ( .A1(n22), .A2(n11), .ZN(n46) );
  INV_X1 U30 ( .A(sel[1]), .ZN(n12) );
  INV_X1 U31 ( .A(sel[2]), .ZN(n4) );
  XNOR2_X1 U32 ( .A(n60), .B(sel[2]), .ZN(n9) );
  XOR2_X1 U33 ( .A(n12), .B(n62), .Z(n13) );
  XOR2_X1 U34 ( .A(sel[2]), .B(A[1]), .Z(n14) );
  XOR2_X1 U35 ( .A(sel[2]), .B(A[2]), .Z(n15) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[1]), .Z(n16) );
  XOR2_X1 U37 ( .A(sel[2]), .B(A[3]), .Z(n17) );
  XOR2_X1 U38 ( .A(sel[1]), .B(A[2]), .Z(n18) );
  XOR2_X1 U39 ( .A(sel[2]), .B(A[4]), .Z(n19) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[3]), .Z(n20) );
  XOR2_X1 U41 ( .A(sel[2]), .B(A[5]), .Z(n21) );
  XOR2_X1 U42 ( .A(sel[1]), .B(A[4]), .Z(n22) );
  XOR2_X1 U43 ( .A(sel[2]), .B(A[6]), .Z(n23) );
  XOR2_X1 U44 ( .A(sel[1]), .B(A[5]), .Z(n24) );
  XOR2_X1 U45 ( .A(sel[2]), .B(A[7]), .Z(n25) );
  XOR2_X1 U46 ( .A(sel[1]), .B(A[6]), .Z(n26) );
  XOR2_X1 U47 ( .A(sel[2]), .B(A[8]), .Z(n27) );
  XOR2_X1 U48 ( .A(sel[1]), .B(A[7]), .Z(n28) );
  XOR2_X1 U49 ( .A(sel[2]), .B(A[9]), .Z(n29) );
  XOR2_X1 U50 ( .A(sel[1]), .B(A[8]), .Z(n30) );
  XOR2_X1 U51 ( .A(sel[2]), .B(A[10]), .Z(n31) );
  XOR2_X1 U52 ( .A(sel[1]), .B(A[9]), .Z(n32) );
  XOR2_X1 U53 ( .A(sel[2]), .B(A[11]), .Z(n33) );
  XOR2_X1 U54 ( .A(sel[1]), .B(A[10]), .Z(n34) );
  XOR2_X1 U55 ( .A(sel[2]), .B(A[12]), .Z(n35) );
  XOR2_X1 U56 ( .A(sel[1]), .B(A[11]), .Z(n36) );
  XOR2_X1 U57 ( .A(sel[2]), .B(A[13]), .Z(n37) );
  XOR2_X1 U58 ( .A(sel[1]), .B(A[12]), .Z(n38) );
  XOR2_X1 U59 ( .A(sel[2]), .B(A[14]), .Z(n39) );
  XOR2_X1 U60 ( .A(sel[1]), .B(A[13]), .Z(n40) );
  XOR2_X1 U61 ( .A(sel[1]), .B(A[14]), .Z(n41) );
  MUX2_X1 U62 ( .A(n42), .B(n14), .S(n8), .Z(B[15]) );
  MUX2_X1 U63 ( .A(n43), .B(n15), .S(n7), .Z(B[16]) );
  MUX2_X1 U64 ( .A(n44), .B(n17), .S(n1), .Z(B[17]) );
  MUX2_X1 U65 ( .A(n45), .B(n19), .S(n8), .Z(B[18]) );
  MUX2_X1 U66 ( .A(n46), .B(n21), .S(n7), .Z(B[19]) );
  MUX2_X1 U67 ( .A(n47), .B(n23), .S(n1), .Z(B[20]) );
  MUX2_X1 U68 ( .A(n48), .B(n25), .S(n8), .Z(B[21]) );
  MUX2_X1 U69 ( .A(n49), .B(n27), .S(n7), .Z(B[22]) );
  MUX2_X1 U70 ( .A(n50), .B(n29), .S(n7), .Z(B[23]) );
  MUX2_X1 U71 ( .A(n51), .B(n31), .S(n1), .Z(B[24]) );
  MUX2_X1 U72 ( .A(n52), .B(n33), .S(n8), .Z(B[25]) );
  MUX2_X1 U73 ( .A(n53), .B(n35), .S(n7), .Z(B[26]) );
  MUX2_X1 U74 ( .A(n54), .B(n37), .S(n1), .Z(B[27]) );
  MUX2_X1 U75 ( .A(n55), .B(n39), .S(n8), .Z(B[28]) );
  MUX2_X1 U76 ( .A(n56), .B(n9), .S(n1), .Z(B[29]) );
  MUX2_X1 U77 ( .A(n10), .B(n58), .S(sel[1]), .Z(n59) );
  OAI21_X1 U78 ( .B1(sel[2]), .B2(n60), .A(sel[0]), .ZN(n57) );
  AOI22_X1 U79 ( .A1(sel[2]), .A2(n60), .B1(sel[0]), .B2(n9), .ZN(n10) );
  INV_X1 U80 ( .A(A[15]), .ZN(n60) );
  AOI21_X1 U81 ( .B1(sel[1]), .B2(sel[0]), .A(n4), .ZN(n63) );
  INV_X1 U82 ( .A(A[0]), .ZN(n62) );
endmodule


module MUX_SHIFT_NB16_N_sh12_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_11, n2, n3, n5, n6, n1, n4, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, \B[0] , n61, n62, n63;
  assign B[31] = B[28];
  assign B[30] = B[28];
  assign B[29] = B[28];
  assign AS = \B[0] ;
  assign B[11] = \B[0] ;
  assign B[10] = \B[0] ;
  assign B[9] = \B[0] ;
  assign B[8] = \B[0] ;
  assign B[7] = \B[0] ;
  assign B[6] = \B[0] ;
  assign B[5] = \B[0] ;
  assign B[4] = \B[0] ;
  assign B[3] = \B[0] ;
  assign B[2] = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  CLKBUF_X3 U3 ( .A(B_11), .Z(\B[0] ) );
  XNOR2_X2 U4 ( .A(n9), .B(sel[0]), .ZN(n4) );
  BUF_X1 U5 ( .A(n61), .Z(n58) );
  BUF_X1 U6 ( .A(n61), .Z(n57) );
  XNOR2_X1 U7 ( .A(n59), .B(n58), .ZN(n1) );
  NOR2_X1 U8 ( .A1(n8), .A2(n10), .ZN(n39) );
  INV_X1 U9 ( .A(A[15]), .ZN(n59) );
  INV_X1 U10 ( .A(n2), .ZN(B[12]) );
  AOI22_X1 U11 ( .A1(n3), .A2(\B[0] ), .B1(n62), .B2(n5), .ZN(n2) );
  INV_X1 U12 ( .A(n3), .ZN(n5) );
  NAND2_X1 U13 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  INV_X1 U14 ( .A(n56), .ZN(B[28]) );
  NAND2_X1 U15 ( .A1(n1), .A2(n54), .ZN(n55) );
  NOR2_X1 U16 ( .A1(n35), .A2(n8), .ZN(n51) );
  NOR2_X1 U17 ( .A1(n13), .A2(n8), .ZN(n40) );
  NOR2_X1 U18 ( .A1(n37), .A2(n8), .ZN(n52) );
  NOR2_X1 U19 ( .A1(n19), .A2(n8), .ZN(n43) );
  NOR2_X1 U20 ( .A1(n21), .A2(n8), .ZN(n44) );
  NOR2_X1 U21 ( .A1(n29), .A2(n8), .ZN(n48) );
  NOR2_X1 U22 ( .A1(n27), .A2(n8), .ZN(n47) );
  NOR2_X1 U23 ( .A1(n33), .A2(n8), .ZN(n50) );
  NOR2_X1 U24 ( .A1(n17), .A2(n8), .ZN(n42) );
  NOR2_X1 U25 ( .A1(n25), .A2(n8), .ZN(n46) );
  NOR2_X1 U27 ( .A1(n38), .A2(n8), .ZN(n53) );
  NOR2_X1 U28 ( .A1(n15), .A2(n8), .ZN(n41) );
  NOR2_X1 U29 ( .A1(n23), .A2(n8), .ZN(n45) );
  NOR2_X1 U30 ( .A1(n31), .A2(n8), .ZN(n49) );
  XOR2_X1 U31 ( .A(n9), .B(n63), .Z(n10) );
  XOR2_X1 U32 ( .A(n58), .B(A[1]), .Z(n11) );
  XOR2_X1 U33 ( .A(n57), .B(A[2]), .Z(n12) );
  XOR2_X1 U34 ( .A(sel[1]), .B(A[1]), .Z(n13) );
  XOR2_X1 U35 ( .A(n57), .B(A[3]), .Z(n14) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[2]), .Z(n15) );
  XOR2_X1 U37 ( .A(n57), .B(A[4]), .Z(n16) );
  XOR2_X1 U38 ( .A(sel[1]), .B(A[3]), .Z(n17) );
  XOR2_X1 U39 ( .A(n58), .B(A[5]), .Z(n18) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[4]), .Z(n19) );
  XOR2_X1 U41 ( .A(n58), .B(A[6]), .Z(n20) );
  XOR2_X1 U42 ( .A(sel[1]), .B(A[5]), .Z(n21) );
  XOR2_X1 U43 ( .A(n58), .B(A[7]), .Z(n22) );
  XOR2_X1 U44 ( .A(sel[1]), .B(A[6]), .Z(n23) );
  XOR2_X1 U45 ( .A(n58), .B(A[8]), .Z(n24) );
  XOR2_X1 U46 ( .A(sel[1]), .B(A[7]), .Z(n25) );
  XOR2_X1 U47 ( .A(n58), .B(A[9]), .Z(n26) );
  XOR2_X1 U48 ( .A(sel[1]), .B(A[8]), .Z(n27) );
  XOR2_X1 U49 ( .A(n58), .B(A[10]), .Z(n28) );
  XOR2_X1 U50 ( .A(sel[1]), .B(A[9]), .Z(n29) );
  XOR2_X1 U51 ( .A(n58), .B(A[11]), .Z(n30) );
  XOR2_X1 U52 ( .A(sel[1]), .B(A[10]), .Z(n31) );
  XOR2_X1 U53 ( .A(n58), .B(A[12]), .Z(n32) );
  XOR2_X1 U54 ( .A(sel[1]), .B(A[11]), .Z(n33) );
  XOR2_X1 U55 ( .A(n58), .B(A[13]), .Z(n34) );
  XOR2_X1 U56 ( .A(sel[1]), .B(A[12]), .Z(n35) );
  XOR2_X1 U57 ( .A(n58), .B(A[14]), .Z(n36) );
  XOR2_X1 U58 ( .A(sel[1]), .B(A[13]), .Z(n37) );
  XOR2_X1 U59 ( .A(sel[1]), .B(A[14]), .Z(n38) );
  MUX2_X1 U60 ( .A(n39), .B(n11), .S(n4), .Z(B[13]) );
  MUX2_X1 U61 ( .A(n40), .B(n12), .S(n4), .Z(B[14]) );
  MUX2_X1 U62 ( .A(n41), .B(n14), .S(n4), .Z(B[15]) );
  MUX2_X1 U63 ( .A(n42), .B(n16), .S(n4), .Z(B[16]) );
  MUX2_X1 U64 ( .A(n43), .B(n18), .S(n4), .Z(B[17]) );
  MUX2_X1 U65 ( .A(n44), .B(n20), .S(n4), .Z(B[18]) );
  MUX2_X1 U66 ( .A(n45), .B(n22), .S(n4), .Z(B[19]) );
  MUX2_X1 U67 ( .A(n46), .B(n24), .S(n4), .Z(B[20]) );
  MUX2_X1 U68 ( .A(n47), .B(n26), .S(n4), .Z(B[21]) );
  MUX2_X1 U69 ( .A(n48), .B(n28), .S(n4), .Z(B[22]) );
  MUX2_X1 U70 ( .A(n49), .B(n30), .S(n4), .Z(B[23]) );
  MUX2_X1 U71 ( .A(n50), .B(n32), .S(n4), .Z(B[24]) );
  MUX2_X1 U72 ( .A(n51), .B(n34), .S(n4), .Z(B[25]) );
  MUX2_X1 U73 ( .A(n52), .B(n36), .S(n4), .Z(B[26]) );
  MUX2_X1 U74 ( .A(n53), .B(n1), .S(n4), .Z(B[27]) );
  MUX2_X1 U75 ( .A(n7), .B(n55), .S(sel[1]), .Z(n56) );
  XOR2_X2 U76 ( .A(n9), .B(n58), .Z(n8) );
  INV_X1 U77 ( .A(sel[1]), .ZN(n9) );
  OAI21_X1 U78 ( .B1(n58), .B2(n59), .A(sel[0]), .ZN(n54) );
  AOI22_X1 U79 ( .A1(n58), .A2(n59), .B1(sel[0]), .B2(n1), .ZN(n7) );
  INV_X1 U80 ( .A(sel[2]), .ZN(n62) );
  AOI21_X1 U81 ( .B1(sel[1]), .B2(sel[0]), .A(n62), .ZN(B_11) );
  INV_X1 U82 ( .A(n62), .ZN(n61) );
  INV_X1 U83 ( .A(A[0]), .ZN(n63) );
endmodule


module MUX_SHIFT_NB16_N_sh10_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_9, n2, n3, n5, n6, n1, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, \B[0] , n61, n62;
  assign B[31] = B[26];
  assign B[30] = B[26];
  assign B[29] = B[26];
  assign B[28] = B[26];
  assign B[27] = B[26];
  assign AS = \B[0] ;
  assign B[9] = \B[0] ;
  assign B[8] = \B[0] ;
  assign B[7] = \B[0] ;
  assign B[6] = \B[0] ;
  assign B[5] = \B[0] ;
  assign B[4] = \B[0] ;
  assign B[3] = \B[0] ;
  assign B[2] = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  CLKBUF_X3 U3 ( .A(B_9), .Z(\B[0] ) );
  XNOR2_X2 U4 ( .A(n9), .B(sel[0]), .ZN(n4) );
  BUF_X1 U5 ( .A(sel[2]), .Z(n58) );
  BUF_X1 U6 ( .A(sel[2]), .Z(n57) );
  XNOR2_X1 U7 ( .A(n59), .B(n58), .ZN(n1) );
  NOR2_X1 U8 ( .A1(n8), .A2(n10), .ZN(n39) );
  INV_X1 U9 ( .A(n2), .ZN(B[10]) );
  AOI22_X1 U10 ( .A1(n3), .A2(\B[0] ), .B1(n61), .B2(n5), .ZN(n2) );
  INV_X1 U11 ( .A(n3), .ZN(n5) );
  NAND2_X1 U12 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  OAI21_X1 U13 ( .B1(n58), .B2(n59), .A(sel[0]), .ZN(n54) );
  NAND2_X1 U14 ( .A1(n1), .A2(n54), .ZN(n55) );
  AOI22_X1 U15 ( .A1(n58), .A2(n59), .B1(sel[0]), .B2(n1), .ZN(n7) );
  NOR2_X1 U16 ( .A1(n38), .A2(n8), .ZN(n53) );
  NOR2_X1 U17 ( .A1(n15), .A2(n8), .ZN(n41) );
  NOR2_X1 U18 ( .A1(n23), .A2(n8), .ZN(n45) );
  NOR2_X1 U19 ( .A1(n17), .A2(n8), .ZN(n42) );
  NOR2_X1 U20 ( .A1(n25), .A2(n8), .ZN(n46) );
  NOR2_X1 U21 ( .A1(n33), .A2(n8), .ZN(n50) );
  NOR2_X1 U22 ( .A1(n31), .A2(n8), .ZN(n49) );
  NOR2_X1 U23 ( .A1(n37), .A2(n8), .ZN(n52) );
  NOR2_X1 U24 ( .A1(n13), .A2(n8), .ZN(n40) );
  NOR2_X1 U25 ( .A1(n21), .A2(n8), .ZN(n44) );
  NOR2_X1 U27 ( .A1(n29), .A2(n8), .ZN(n48) );
  NOR2_X1 U28 ( .A1(n19), .A2(n8), .ZN(n43) );
  NOR2_X1 U29 ( .A1(n27), .A2(n8), .ZN(n47) );
  NOR2_X1 U30 ( .A1(n35), .A2(n8), .ZN(n51) );
  XOR2_X1 U31 ( .A(n9), .B(n62), .Z(n10) );
  XOR2_X1 U32 ( .A(n58), .B(A[1]), .Z(n11) );
  XOR2_X1 U33 ( .A(n57), .B(A[2]), .Z(n12) );
  XOR2_X1 U34 ( .A(sel[1]), .B(A[1]), .Z(n13) );
  XOR2_X1 U35 ( .A(n57), .B(A[3]), .Z(n14) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[2]), .Z(n15) );
  XOR2_X1 U37 ( .A(n57), .B(A[4]), .Z(n16) );
  XOR2_X1 U38 ( .A(sel[1]), .B(A[3]), .Z(n17) );
  XOR2_X1 U39 ( .A(n58), .B(A[5]), .Z(n18) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[4]), .Z(n19) );
  XOR2_X1 U41 ( .A(n58), .B(A[6]), .Z(n20) );
  XOR2_X1 U42 ( .A(sel[1]), .B(A[5]), .Z(n21) );
  XOR2_X1 U43 ( .A(n58), .B(A[7]), .Z(n22) );
  XOR2_X1 U44 ( .A(sel[1]), .B(A[6]), .Z(n23) );
  XOR2_X1 U45 ( .A(n58), .B(A[8]), .Z(n24) );
  XOR2_X1 U46 ( .A(sel[1]), .B(A[7]), .Z(n25) );
  XOR2_X1 U47 ( .A(n58), .B(A[9]), .Z(n26) );
  XOR2_X1 U48 ( .A(sel[1]), .B(A[8]), .Z(n27) );
  XOR2_X1 U49 ( .A(n58), .B(A[10]), .Z(n28) );
  XOR2_X1 U50 ( .A(sel[1]), .B(A[9]), .Z(n29) );
  XOR2_X1 U51 ( .A(n58), .B(A[11]), .Z(n30) );
  XOR2_X1 U52 ( .A(sel[1]), .B(A[10]), .Z(n31) );
  XOR2_X1 U53 ( .A(n58), .B(A[12]), .Z(n32) );
  XOR2_X1 U54 ( .A(sel[1]), .B(A[11]), .Z(n33) );
  XOR2_X1 U55 ( .A(n58), .B(A[13]), .Z(n34) );
  XOR2_X1 U56 ( .A(sel[1]), .B(A[12]), .Z(n35) );
  XOR2_X1 U57 ( .A(n58), .B(A[14]), .Z(n36) );
  XOR2_X1 U58 ( .A(sel[1]), .B(A[13]), .Z(n37) );
  XOR2_X1 U59 ( .A(sel[1]), .B(A[14]), .Z(n38) );
  MUX2_X1 U60 ( .A(n39), .B(n11), .S(n4), .Z(B[11]) );
  MUX2_X1 U61 ( .A(n40), .B(n12), .S(n4), .Z(B[12]) );
  MUX2_X1 U62 ( .A(n41), .B(n14), .S(n4), .Z(B[13]) );
  MUX2_X1 U63 ( .A(n42), .B(n16), .S(n4), .Z(B[14]) );
  MUX2_X1 U64 ( .A(n43), .B(n18), .S(n4), .Z(B[15]) );
  MUX2_X1 U65 ( .A(n44), .B(n20), .S(n4), .Z(B[16]) );
  MUX2_X1 U66 ( .A(n45), .B(n22), .S(n4), .Z(B[17]) );
  MUX2_X1 U67 ( .A(n46), .B(n24), .S(n4), .Z(B[18]) );
  MUX2_X1 U68 ( .A(n47), .B(n26), .S(n4), .Z(B[19]) );
  MUX2_X1 U69 ( .A(n48), .B(n28), .S(n4), .Z(B[20]) );
  MUX2_X1 U70 ( .A(n49), .B(n30), .S(n4), .Z(B[21]) );
  MUX2_X1 U71 ( .A(n50), .B(n32), .S(n4), .Z(B[22]) );
  MUX2_X1 U72 ( .A(n51), .B(n34), .S(n4), .Z(B[23]) );
  MUX2_X1 U73 ( .A(n52), .B(n36), .S(n4), .Z(B[24]) );
  MUX2_X1 U74 ( .A(n53), .B(n1), .S(n4), .Z(B[25]) );
  MUX2_X1 U75 ( .A(n7), .B(n55), .S(sel[1]), .Z(n56) );
  INV_X2 U76 ( .A(n56), .ZN(B[26]) );
  XOR2_X2 U77 ( .A(n9), .B(n58), .Z(n8) );
  INV_X1 U78 ( .A(sel[1]), .ZN(n9) );
  INV_X1 U79 ( .A(A[15]), .ZN(n59) );
  INV_X1 U80 ( .A(sel[2]), .ZN(n61) );
  AOI21_X1 U81 ( .B1(sel[0]), .B2(sel[1]), .A(n61), .ZN(B_9) );
  INV_X1 U82 ( .A(A[0]), .ZN(n62) );
endmodule


module MUX_SHIFT_NB16_N_sh8_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_7, n2, n3, n5, n6, n1, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, \B[0] , n61, n62;
  assign B[31] = B[24];
  assign B[30] = B[24];
  assign B[29] = B[24];
  assign B[28] = B[24];
  assign B[27] = B[24];
  assign B[26] = B[24];
  assign B[25] = B[24];
  assign AS = \B[0] ;
  assign B[7] = \B[0] ;
  assign B[6] = \B[0] ;
  assign B[5] = \B[0] ;
  assign B[4] = \B[0] ;
  assign B[3] = \B[0] ;
  assign B[2] = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  XNOR2_X2 U3 ( .A(n9), .B(sel[0]), .ZN(n4) );
  BUF_X2 U4 ( .A(B_7), .Z(\B[0] ) );
  BUF_X1 U5 ( .A(sel[2]), .Z(n58) );
  BUF_X1 U6 ( .A(sel[2]), .Z(n57) );
  XNOR2_X1 U7 ( .A(n59), .B(n58), .ZN(n1) );
  NOR2_X1 U8 ( .A1(n8), .A2(n10), .ZN(n39) );
  INV_X1 U9 ( .A(n2), .ZN(B[8]) );
  AOI22_X1 U10 ( .A1(n3), .A2(\B[0] ), .B1(n61), .B2(n5), .ZN(n2) );
  INV_X1 U11 ( .A(n3), .ZN(n5) );
  NAND2_X1 U12 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  INV_X1 U13 ( .A(sel[2]), .ZN(n61) );
  NAND2_X1 U14 ( .A1(n1), .A2(n54), .ZN(n55) );
  AOI22_X1 U15 ( .A1(n58), .A2(n59), .B1(sel[0]), .B2(n1), .ZN(n7) );
  AOI21_X1 U16 ( .B1(sel[1]), .B2(sel[0]), .A(n61), .ZN(B_7) );
  NOR2_X1 U17 ( .A1(n13), .A2(n8), .ZN(n40) );
  NOR2_X1 U18 ( .A1(n19), .A2(n8), .ZN(n43) );
  NOR2_X1 U19 ( .A1(n27), .A2(n8), .ZN(n47) );
  NOR2_X1 U20 ( .A1(n21), .A2(n8), .ZN(n44) );
  NOR2_X1 U21 ( .A1(n29), .A2(n8), .ZN(n48) );
  NOR2_X1 U22 ( .A1(n37), .A2(n8), .ZN(n52) );
  NOR2_X1 U23 ( .A1(n35), .A2(n8), .ZN(n51) );
  NOR2_X1 U24 ( .A1(n17), .A2(n8), .ZN(n42) );
  NOR2_X1 U25 ( .A1(n25), .A2(n8), .ZN(n46) );
  NOR2_X1 U27 ( .A1(n33), .A2(n8), .ZN(n50) );
  NOR2_X1 U28 ( .A1(n15), .A2(n8), .ZN(n41) );
  NOR2_X1 U29 ( .A1(n23), .A2(n8), .ZN(n45) );
  NOR2_X1 U30 ( .A1(n31), .A2(n8), .ZN(n49) );
  NOR2_X1 U31 ( .A1(n38), .A2(n8), .ZN(n53) );
  OAI21_X1 U32 ( .B1(n58), .B2(n59), .A(sel[0]), .ZN(n54) );
  INV_X1 U33 ( .A(sel[1]), .ZN(n9) );
  XOR2_X1 U34 ( .A(n9), .B(n62), .Z(n10) );
  XOR2_X1 U35 ( .A(n58), .B(A[1]), .Z(n11) );
  XOR2_X1 U36 ( .A(n57), .B(A[2]), .Z(n12) );
  XOR2_X1 U37 ( .A(sel[1]), .B(A[1]), .Z(n13) );
  XOR2_X1 U38 ( .A(n57), .B(A[3]), .Z(n14) );
  XOR2_X1 U39 ( .A(sel[1]), .B(A[2]), .Z(n15) );
  XOR2_X1 U40 ( .A(n57), .B(A[4]), .Z(n16) );
  XOR2_X1 U41 ( .A(sel[1]), .B(A[3]), .Z(n17) );
  XOR2_X1 U42 ( .A(n58), .B(A[5]), .Z(n18) );
  XOR2_X1 U43 ( .A(sel[1]), .B(A[4]), .Z(n19) );
  XOR2_X1 U44 ( .A(n58), .B(A[6]), .Z(n20) );
  XOR2_X1 U45 ( .A(sel[1]), .B(A[5]), .Z(n21) );
  XOR2_X1 U46 ( .A(n58), .B(A[7]), .Z(n22) );
  XOR2_X1 U47 ( .A(sel[1]), .B(A[6]), .Z(n23) );
  XOR2_X1 U48 ( .A(n58), .B(A[8]), .Z(n24) );
  XOR2_X1 U49 ( .A(sel[1]), .B(A[7]), .Z(n25) );
  XOR2_X1 U50 ( .A(n58), .B(A[9]), .Z(n26) );
  XOR2_X1 U51 ( .A(sel[1]), .B(A[8]), .Z(n27) );
  XOR2_X1 U52 ( .A(n58), .B(A[10]), .Z(n28) );
  XOR2_X1 U53 ( .A(sel[1]), .B(A[9]), .Z(n29) );
  XOR2_X1 U54 ( .A(n58), .B(A[11]), .Z(n30) );
  XOR2_X1 U55 ( .A(sel[1]), .B(A[10]), .Z(n31) );
  XOR2_X1 U56 ( .A(n58), .B(A[12]), .Z(n32) );
  XOR2_X1 U57 ( .A(sel[1]), .B(A[11]), .Z(n33) );
  XOR2_X1 U58 ( .A(n58), .B(A[13]), .Z(n34) );
  XOR2_X1 U59 ( .A(sel[1]), .B(A[12]), .Z(n35) );
  XOR2_X1 U60 ( .A(n58), .B(A[14]), .Z(n36) );
  XOR2_X1 U61 ( .A(sel[1]), .B(A[13]), .Z(n37) );
  XOR2_X1 U62 ( .A(sel[1]), .B(A[14]), .Z(n38) );
  MUX2_X1 U63 ( .A(n39), .B(n11), .S(n4), .Z(B[9]) );
  MUX2_X1 U64 ( .A(n40), .B(n12), .S(n4), .Z(B[10]) );
  MUX2_X1 U65 ( .A(n41), .B(n14), .S(n4), .Z(B[11]) );
  MUX2_X1 U66 ( .A(n42), .B(n16), .S(n4), .Z(B[12]) );
  MUX2_X1 U67 ( .A(n43), .B(n18), .S(n4), .Z(B[13]) );
  MUX2_X1 U68 ( .A(n44), .B(n20), .S(n4), .Z(B[14]) );
  MUX2_X1 U69 ( .A(n45), .B(n22), .S(n4), .Z(B[15]) );
  MUX2_X1 U70 ( .A(n46), .B(n24), .S(n4), .Z(B[16]) );
  MUX2_X1 U71 ( .A(n47), .B(n26), .S(n4), .Z(B[17]) );
  MUX2_X1 U72 ( .A(n48), .B(n28), .S(n4), .Z(B[18]) );
  MUX2_X1 U73 ( .A(n49), .B(n30), .S(n4), .Z(B[19]) );
  MUX2_X1 U74 ( .A(n50), .B(n32), .S(n4), .Z(B[20]) );
  MUX2_X1 U75 ( .A(n51), .B(n34), .S(n4), .Z(B[21]) );
  MUX2_X1 U76 ( .A(n52), .B(n36), .S(n4), .Z(B[22]) );
  MUX2_X1 U77 ( .A(n53), .B(n1), .S(n4), .Z(B[23]) );
  MUX2_X1 U78 ( .A(n7), .B(n55), .S(sel[1]), .Z(n56) );
  INV_X2 U79 ( .A(n56), .ZN(B[24]) );
  XOR2_X2 U80 ( .A(n9), .B(n58), .Z(n8) );
  INV_X1 U81 ( .A(A[15]), .ZN(n59) );
  INV_X1 U82 ( .A(A[0]), .ZN(n62) );
endmodule


module MUX_SHIFT_NB16_N_sh6_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_5, n2, n3, n5, n6, n1, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, \B[0] , n61, n62;
  assign B[31] = B[22];
  assign B[30] = B[22];
  assign B[29] = B[22];
  assign B[28] = B[22];
  assign B[27] = B[22];
  assign B[26] = B[22];
  assign B[25] = B[22];
  assign B[24] = B[22];
  assign B[23] = B[22];
  assign AS = \B[0] ;
  assign B[5] = \B[0] ;
  assign B[4] = \B[0] ;
  assign B[3] = \B[0] ;
  assign B[2] = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  BUF_X2 U3 ( .A(n7), .Z(B[22]) );
  XNOR2_X2 U4 ( .A(n10), .B(sel[0]), .ZN(n4) );
  BUF_X1 U5 ( .A(sel[2]), .Z(n58) );
  XNOR2_X1 U6 ( .A(n59), .B(n58), .ZN(n1) );
  NOR2_X1 U7 ( .A1(n9), .A2(n11), .ZN(n40) );
  INV_X1 U8 ( .A(n2), .ZN(B[6]) );
  AOI22_X1 U9 ( .A1(n3), .A2(\B[0] ), .B1(n61), .B2(n5), .ZN(n2) );
  INV_X1 U10 ( .A(n3), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  BUF_X2 U12 ( .A(B_5), .Z(\B[0] ) );
  NOR2_X1 U13 ( .A1(n16), .A2(n9), .ZN(n42) );
  NOR2_X1 U14 ( .A1(n18), .A2(n9), .ZN(n43) );
  NOR2_X1 U15 ( .A1(n24), .A2(n9), .ZN(n46) );
  NOR2_X1 U16 ( .A1(n32), .A2(n9), .ZN(n50) );
  NOR2_X1 U17 ( .A1(n26), .A2(n9), .ZN(n47) );
  NOR2_X1 U18 ( .A1(n34), .A2(n9), .ZN(n51) );
  NOR2_X1 U19 ( .A1(n39), .A2(n9), .ZN(n54) );
  NOR2_X1 U20 ( .A1(n14), .A2(n9), .ZN(n41) );
  NOR2_X1 U21 ( .A1(n22), .A2(n9), .ZN(n45) );
  NOR2_X1 U22 ( .A1(n30), .A2(n9), .ZN(n49) );
  NOR2_X1 U23 ( .A1(n38), .A2(n9), .ZN(n53) );
  NOR2_X1 U24 ( .A1(n20), .A2(n9), .ZN(n44) );
  NOR2_X1 U25 ( .A1(n28), .A2(n9), .ZN(n48) );
  NOR2_X1 U27 ( .A1(n36), .A2(n9), .ZN(n52) );
  INV_X1 U28 ( .A(sel[2]), .ZN(n61) );
  INV_X1 U29 ( .A(n57), .ZN(n7) );
  NAND2_X1 U30 ( .A1(n1), .A2(n55), .ZN(n56) );
  XOR2_X1 U31 ( .A(n10), .B(n62), .Z(n11) );
  XOR2_X1 U32 ( .A(n58), .B(A[1]), .Z(n12) );
  XOR2_X1 U33 ( .A(n58), .B(A[2]), .Z(n13) );
  XOR2_X1 U34 ( .A(sel[1]), .B(A[1]), .Z(n14) );
  XOR2_X1 U35 ( .A(n58), .B(A[3]), .Z(n15) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[2]), .Z(n16) );
  XOR2_X1 U37 ( .A(n58), .B(A[4]), .Z(n17) );
  XOR2_X1 U38 ( .A(sel[1]), .B(A[3]), .Z(n18) );
  XOR2_X1 U39 ( .A(n58), .B(A[5]), .Z(n19) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[4]), .Z(n20) );
  XOR2_X1 U41 ( .A(n58), .B(A[6]), .Z(n21) );
  XOR2_X1 U42 ( .A(sel[1]), .B(A[5]), .Z(n22) );
  XOR2_X1 U43 ( .A(n58), .B(A[7]), .Z(n23) );
  XOR2_X1 U44 ( .A(sel[1]), .B(A[6]), .Z(n24) );
  XOR2_X1 U45 ( .A(n58), .B(A[8]), .Z(n25) );
  XOR2_X1 U46 ( .A(sel[1]), .B(A[7]), .Z(n26) );
  XOR2_X1 U47 ( .A(n58), .B(A[9]), .Z(n27) );
  XOR2_X1 U48 ( .A(sel[1]), .B(A[8]), .Z(n28) );
  XOR2_X1 U49 ( .A(n58), .B(A[10]), .Z(n29) );
  XOR2_X1 U50 ( .A(sel[1]), .B(A[9]), .Z(n30) );
  XOR2_X1 U51 ( .A(n58), .B(A[11]), .Z(n31) );
  XOR2_X1 U52 ( .A(sel[1]), .B(A[10]), .Z(n32) );
  XOR2_X1 U53 ( .A(n58), .B(A[12]), .Z(n33) );
  XOR2_X1 U54 ( .A(sel[1]), .B(A[11]), .Z(n34) );
  XOR2_X1 U55 ( .A(n58), .B(A[13]), .Z(n35) );
  XOR2_X1 U56 ( .A(sel[1]), .B(A[12]), .Z(n36) );
  XOR2_X1 U57 ( .A(n58), .B(A[14]), .Z(n37) );
  XOR2_X1 U58 ( .A(sel[1]), .B(A[13]), .Z(n38) );
  XOR2_X1 U59 ( .A(sel[1]), .B(A[14]), .Z(n39) );
  MUX2_X1 U60 ( .A(n40), .B(n12), .S(n4), .Z(B[7]) );
  MUX2_X1 U61 ( .A(n41), .B(n13), .S(n4), .Z(B[8]) );
  MUX2_X1 U62 ( .A(n42), .B(n15), .S(n4), .Z(B[9]) );
  MUX2_X1 U63 ( .A(n43), .B(n17), .S(n4), .Z(B[10]) );
  MUX2_X1 U64 ( .A(n44), .B(n19), .S(n4), .Z(B[11]) );
  MUX2_X1 U65 ( .A(n45), .B(n21), .S(n4), .Z(B[12]) );
  MUX2_X1 U66 ( .A(n46), .B(n23), .S(n4), .Z(B[13]) );
  MUX2_X1 U67 ( .A(n47), .B(n25), .S(n4), .Z(B[14]) );
  MUX2_X1 U68 ( .A(n48), .B(n27), .S(n4), .Z(B[15]) );
  MUX2_X1 U69 ( .A(n49), .B(n29), .S(n4), .Z(B[16]) );
  MUX2_X1 U70 ( .A(n50), .B(n31), .S(n4), .Z(B[17]) );
  MUX2_X1 U71 ( .A(n51), .B(n33), .S(n4), .Z(B[18]) );
  MUX2_X1 U72 ( .A(n52), .B(n35), .S(n4), .Z(B[19]) );
  MUX2_X1 U73 ( .A(n53), .B(n37), .S(n4), .Z(B[20]) );
  MUX2_X1 U74 ( .A(n54), .B(n1), .S(n4), .Z(B[21]) );
  MUX2_X1 U75 ( .A(n8), .B(n56), .S(sel[1]), .Z(n57) );
  XOR2_X2 U76 ( .A(n10), .B(n58), .Z(n9) );
  INV_X1 U77 ( .A(sel[1]), .ZN(n10) );
  OAI21_X1 U78 ( .B1(n58), .B2(n59), .A(sel[0]), .ZN(n55) );
  AOI22_X1 U79 ( .A1(n58), .A2(n59), .B1(sel[0]), .B2(n1), .ZN(n8) );
  INV_X1 U80 ( .A(A[15]), .ZN(n59) );
  AOI21_X1 U81 ( .B1(sel[1]), .B2(sel[0]), .A(n61), .ZN(B_5) );
  INV_X1 U82 ( .A(A[0]), .ZN(n62) );
endmodule


module MUX_SHIFT_NB16_N_sh4_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_3, n2, n3, n5, n6, n1, n4, \B[20] , n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, \B[0] , n63, n64;
  assign B[31] = \B[20] ;
  assign B[30] = \B[20] ;
  assign B[29] = \B[20] ;
  assign B[28] = \B[20] ;
  assign B[27] = \B[20] ;
  assign B[26] = \B[20] ;
  assign B[25] = \B[20] ;
  assign B[24] = \B[20] ;
  assign B[23] = \B[20] ;
  assign B[22] = \B[20] ;
  assign B[21] = \B[20] ;
  assign B[20] = \B[20] ;
  assign AS = \B[0] ;
  assign B[3] = \B[0] ;
  assign B[2] = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  INV_X4 U3 ( .A(n56), .ZN(\B[20] ) );
  XNOR2_X2 U4 ( .A(n58), .B(sel[0]), .ZN(n4) );
  BUF_X1 U5 ( .A(B_3), .Z(\B[0] ) );
  INV_X1 U6 ( .A(n58), .ZN(n60) );
  BUF_X1 U7 ( .A(sel[2]), .Z(n57) );
  XNOR2_X1 U8 ( .A(n61), .B(n57), .ZN(n1) );
  NOR2_X1 U9 ( .A1(n19), .A2(n9), .ZN(n43) );
  NOR2_X1 U10 ( .A1(n21), .A2(n9), .ZN(n44) );
  NOR2_X1 U11 ( .A1(n9), .A2(n10), .ZN(n39) );
  NOR2_X1 U12 ( .A1(n27), .A2(n9), .ZN(n47) );
  NOR2_X1 U13 ( .A1(n13), .A2(n9), .ZN(n40) );
  NOR2_X1 U14 ( .A1(n35), .A2(n9), .ZN(n51) );
  NOR2_X1 U15 ( .A1(n29), .A2(n9), .ZN(n48) );
  NOR2_X1 U16 ( .A1(n37), .A2(n9), .ZN(n52) );
  NOR2_X1 U17 ( .A1(n17), .A2(n9), .ZN(n42) );
  NOR2_X1 U18 ( .A1(n25), .A2(n9), .ZN(n46) );
  NOR2_X1 U19 ( .A1(n33), .A2(n9), .ZN(n50) );
  NOR2_X1 U20 ( .A1(n23), .A2(n9), .ZN(n45) );
  NOR2_X1 U21 ( .A1(n15), .A2(n9), .ZN(n41) );
  NOR2_X1 U22 ( .A1(n31), .A2(n9), .ZN(n49) );
  NOR2_X1 U23 ( .A1(n38), .A2(n9), .ZN(n53) );
  INV_X1 U24 ( .A(n2), .ZN(B[4]) );
  AOI22_X1 U25 ( .A1(n3), .A2(\B[0] ), .B1(n63), .B2(n5), .ZN(n2) );
  INV_X1 U27 ( .A(n3), .ZN(n5) );
  NAND2_X1 U28 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  NAND2_X1 U29 ( .A1(n1), .A2(n54), .ZN(n55) );
  XOR2_X1 U30 ( .A(n58), .B(n64), .Z(n10) );
  XOR2_X1 U31 ( .A(n57), .B(A[1]), .Z(n11) );
  XOR2_X1 U32 ( .A(n57), .B(A[2]), .Z(n12) );
  XOR2_X1 U33 ( .A(n60), .B(A[1]), .Z(n13) );
  XOR2_X1 U34 ( .A(n57), .B(A[3]), .Z(n14) );
  XOR2_X1 U35 ( .A(n60), .B(A[2]), .Z(n15) );
  XOR2_X1 U36 ( .A(n57), .B(A[4]), .Z(n16) );
  XOR2_X1 U37 ( .A(n60), .B(A[3]), .Z(n17) );
  XOR2_X1 U38 ( .A(n57), .B(A[5]), .Z(n18) );
  XOR2_X1 U39 ( .A(n60), .B(A[4]), .Z(n19) );
  XOR2_X1 U40 ( .A(n57), .B(A[6]), .Z(n20) );
  XOR2_X1 U41 ( .A(n60), .B(A[5]), .Z(n21) );
  XOR2_X1 U42 ( .A(n57), .B(A[7]), .Z(n22) );
  XOR2_X1 U43 ( .A(n60), .B(A[6]), .Z(n23) );
  XOR2_X1 U44 ( .A(n57), .B(A[8]), .Z(n24) );
  XOR2_X1 U45 ( .A(n60), .B(A[7]), .Z(n25) );
  XOR2_X1 U46 ( .A(n57), .B(A[9]), .Z(n26) );
  XOR2_X1 U47 ( .A(n60), .B(A[8]), .Z(n27) );
  XOR2_X1 U48 ( .A(n57), .B(A[10]), .Z(n28) );
  XOR2_X1 U49 ( .A(n60), .B(A[9]), .Z(n29) );
  XOR2_X1 U50 ( .A(n57), .B(A[11]), .Z(n30) );
  XOR2_X1 U51 ( .A(n60), .B(A[10]), .Z(n31) );
  XOR2_X1 U52 ( .A(n57), .B(A[12]), .Z(n32) );
  XOR2_X1 U53 ( .A(n60), .B(A[11]), .Z(n33) );
  XOR2_X1 U54 ( .A(n57), .B(A[13]), .Z(n34) );
  XOR2_X1 U55 ( .A(n60), .B(A[12]), .Z(n35) );
  XOR2_X1 U56 ( .A(n57), .B(A[14]), .Z(n36) );
  XOR2_X1 U57 ( .A(n59), .B(A[13]), .Z(n37) );
  XOR2_X1 U58 ( .A(n59), .B(A[14]), .Z(n38) );
  MUX2_X1 U59 ( .A(n39), .B(n11), .S(n4), .Z(B[5]) );
  MUX2_X1 U60 ( .A(n40), .B(n12), .S(n4), .Z(B[6]) );
  MUX2_X1 U61 ( .A(n41), .B(n14), .S(n4), .Z(B[7]) );
  MUX2_X1 U62 ( .A(n42), .B(n16), .S(n4), .Z(B[8]) );
  MUX2_X1 U63 ( .A(n43), .B(n18), .S(n4), .Z(B[9]) );
  MUX2_X1 U64 ( .A(n44), .B(n20), .S(n4), .Z(B[10]) );
  MUX2_X1 U65 ( .A(n45), .B(n22), .S(n4), .Z(B[11]) );
  MUX2_X1 U66 ( .A(n46), .B(n24), .S(n4), .Z(B[12]) );
  MUX2_X1 U67 ( .A(n47), .B(n26), .S(n4), .Z(B[13]) );
  MUX2_X1 U68 ( .A(n48), .B(n28), .S(n4), .Z(B[14]) );
  MUX2_X1 U69 ( .A(n49), .B(n30), .S(n4), .Z(B[15]) );
  MUX2_X1 U70 ( .A(n50), .B(n32), .S(n4), .Z(B[16]) );
  MUX2_X1 U71 ( .A(n51), .B(n34), .S(n4), .Z(B[17]) );
  MUX2_X1 U72 ( .A(n52), .B(n36), .S(n4), .Z(B[18]) );
  MUX2_X1 U73 ( .A(n53), .B(n1), .S(n4), .Z(B[19]) );
  MUX2_X1 U74 ( .A(n8), .B(n55), .S(n59), .Z(n56) );
  INV_X1 U75 ( .A(sel[1]), .ZN(n58) );
  INV_X1 U76 ( .A(n58), .ZN(n59) );
  XOR2_X2 U77 ( .A(n58), .B(n57), .Z(n9) );
  OAI21_X1 U78 ( .B1(n57), .B2(n61), .A(sel[0]), .ZN(n54) );
  AOI22_X1 U79 ( .A1(n57), .A2(n61), .B1(sel[0]), .B2(n1), .ZN(n8) );
  INV_X1 U80 ( .A(A[15]), .ZN(n61) );
  AOI21_X1 U81 ( .B1(sel[1]), .B2(sel[0]), .A(n63), .ZN(B_3) );
  INV_X1 U82 ( .A(sel[2]), .ZN(n63) );
  INV_X1 U83 ( .A(A[0]), .ZN(n64) );
endmodule


module MUX_SHIFT_NB16_N_sh2_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_1, n2, n3, n5, n6, n1, n4, \B[0] , n8, \B[18] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64;
  assign AS = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;
  assign B[31] = \B[18] ;
  assign B[30] = \B[18] ;
  assign B[29] = \B[18] ;
  assign B[28] = \B[18] ;
  assign B[27] = \B[18] ;
  assign B[26] = \B[18] ;
  assign B[25] = \B[18] ;
  assign B[24] = \B[18] ;
  assign B[23] = \B[18] ;
  assign B[22] = \B[18] ;
  assign B[21] = \B[18] ;
  assign B[20] = \B[18] ;
  assign B[19] = \B[18] ;
  assign B[18] = \B[18] ;

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  INV_X4 U3 ( .A(n58), .ZN(\B[18] ) );
  XOR2_X1 U4 ( .A(n60), .B(sel[0]), .Z(n1) );
  INV_X1 U5 ( .A(n1), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(B_1), .Z(\B[0] ) );
  AOI21_X1 U7 ( .B1(sel[1]), .B2(sel[0]), .A(n63), .ZN(B_1) );
  INV_X1 U8 ( .A(n60), .ZN(n61) );
  BUF_X1 U9 ( .A(sel[2]), .Z(n59) );
  XNOR2_X1 U10 ( .A(n62), .B(n59), .ZN(n8) );
  NOR2_X1 U11 ( .A1(n25), .A2(n11), .ZN(n47) );
  NOR2_X1 U12 ( .A1(n27), .A2(n11), .ZN(n48) );
  NOR2_X1 U13 ( .A1(n17), .A2(n11), .ZN(n43) );
  NOR2_X1 U14 ( .A1(n33), .A2(n11), .ZN(n51) );
  NOR2_X1 U15 ( .A1(n19), .A2(n11), .ZN(n44) );
  NOR2_X1 U16 ( .A1(n40), .A2(n11), .ZN(n55) );
  NOR2_X1 U17 ( .A1(n35), .A2(n11), .ZN(n52) );
  NOR2_X1 U18 ( .A1(n23), .A2(n11), .ZN(n46) );
  NOR2_X1 U19 ( .A1(n15), .A2(n11), .ZN(n42) );
  NOR2_X1 U20 ( .A1(n31), .A2(n11), .ZN(n50) );
  NOR2_X1 U21 ( .A1(n39), .A2(n11), .ZN(n54) );
  INV_X1 U22 ( .A(n2), .ZN(B[2]) );
  AOI22_X1 U23 ( .A1(n3), .A2(\B[0] ), .B1(n63), .B2(n5), .ZN(n2) );
  INV_X1 U24 ( .A(n3), .ZN(n5) );
  NAND2_X1 U25 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  NOR2_X1 U27 ( .A1(n29), .A2(n11), .ZN(n49) );
  NOR2_X1 U28 ( .A1(n11), .A2(n12), .ZN(n41) );
  NOR2_X1 U29 ( .A1(n21), .A2(n11), .ZN(n45) );
  NOR2_X1 U30 ( .A1(n37), .A2(n11), .ZN(n53) );
  NAND2_X1 U31 ( .A1(n8), .A2(n56), .ZN(n57) );
  XOR2_X1 U32 ( .A(n60), .B(n64), .Z(n12) );
  XOR2_X1 U33 ( .A(n59), .B(A[1]), .Z(n13) );
  XOR2_X1 U34 ( .A(n59), .B(A[2]), .Z(n14) );
  XOR2_X1 U35 ( .A(n61), .B(A[1]), .Z(n15) );
  XOR2_X1 U36 ( .A(n59), .B(A[3]), .Z(n16) );
  XOR2_X1 U37 ( .A(n61), .B(A[2]), .Z(n17) );
  XOR2_X1 U38 ( .A(n59), .B(A[4]), .Z(n18) );
  XOR2_X1 U39 ( .A(n61), .B(A[3]), .Z(n19) );
  XOR2_X1 U40 ( .A(n59), .B(A[5]), .Z(n20) );
  XOR2_X1 U41 ( .A(n61), .B(A[4]), .Z(n21) );
  XOR2_X1 U42 ( .A(n59), .B(A[6]), .Z(n22) );
  XOR2_X1 U43 ( .A(n61), .B(A[5]), .Z(n23) );
  XOR2_X1 U44 ( .A(n59), .B(A[7]), .Z(n24) );
  XOR2_X1 U45 ( .A(n61), .B(A[6]), .Z(n25) );
  XOR2_X1 U46 ( .A(n59), .B(A[8]), .Z(n26) );
  XOR2_X1 U47 ( .A(n61), .B(A[7]), .Z(n27) );
  XOR2_X1 U48 ( .A(n59), .B(A[9]), .Z(n28) );
  XOR2_X1 U49 ( .A(n61), .B(A[8]), .Z(n29) );
  XOR2_X1 U50 ( .A(n59), .B(A[10]), .Z(n30) );
  XOR2_X1 U51 ( .A(n61), .B(A[9]), .Z(n31) );
  XOR2_X1 U52 ( .A(n59), .B(A[11]), .Z(n32) );
  XOR2_X1 U53 ( .A(n61), .B(A[10]), .Z(n33) );
  XOR2_X1 U54 ( .A(n59), .B(A[12]), .Z(n34) );
  XOR2_X1 U55 ( .A(n61), .B(A[11]), .Z(n35) );
  XOR2_X1 U56 ( .A(n59), .B(A[13]), .Z(n36) );
  XOR2_X1 U57 ( .A(n61), .B(A[12]), .Z(n37) );
  XOR2_X1 U58 ( .A(n59), .B(A[14]), .Z(n38) );
  XOR2_X1 U59 ( .A(sel[1]), .B(A[13]), .Z(n39) );
  XOR2_X1 U60 ( .A(sel[1]), .B(A[14]), .Z(n40) );
  MUX2_X1 U61 ( .A(n41), .B(n13), .S(n4), .Z(B[3]) );
  MUX2_X1 U62 ( .A(n42), .B(n14), .S(n4), .Z(B[4]) );
  MUX2_X1 U63 ( .A(n43), .B(n16), .S(n4), .Z(B[5]) );
  MUX2_X1 U64 ( .A(n44), .B(n18), .S(n4), .Z(B[6]) );
  MUX2_X1 U65 ( .A(n45), .B(n20), .S(n4), .Z(B[7]) );
  MUX2_X1 U66 ( .A(n46), .B(n22), .S(n4), .Z(B[8]) );
  MUX2_X1 U67 ( .A(n47), .B(n24), .S(n4), .Z(B[9]) );
  MUX2_X1 U68 ( .A(n48), .B(n26), .S(n4), .Z(B[10]) );
  MUX2_X1 U69 ( .A(n49), .B(n28), .S(n4), .Z(B[11]) );
  MUX2_X1 U70 ( .A(n50), .B(n30), .S(n4), .Z(B[12]) );
  MUX2_X1 U71 ( .A(n51), .B(n32), .S(n4), .Z(B[13]) );
  MUX2_X1 U72 ( .A(n52), .B(n34), .S(n4), .Z(B[14]) );
  MUX2_X1 U73 ( .A(n53), .B(n36), .S(n4), .Z(B[15]) );
  MUX2_X1 U74 ( .A(n54), .B(n38), .S(n4), .Z(B[16]) );
  MUX2_X1 U75 ( .A(n55), .B(n8), .S(n4), .Z(B[17]) );
  MUX2_X1 U76 ( .A(n10), .B(n57), .S(sel[1]), .Z(n58) );
  INV_X1 U77 ( .A(sel[1]), .ZN(n60) );
  XOR2_X2 U78 ( .A(n60), .B(n59), .Z(n11) );
  OAI21_X1 U79 ( .B1(n59), .B2(n62), .A(sel[0]), .ZN(n56) );
  AOI22_X1 U80 ( .A1(n59), .A2(n62), .B1(sel[0]), .B2(n8), .ZN(n10) );
  INV_X1 U81 ( .A(A[15]), .ZN(n62) );
  INV_X1 U82 ( .A(sel[2]), .ZN(n63) );
  INV_X1 U83 ( .A(A[0]), .ZN(n64) );
endmodule


module MUX_SHIFT_NB16_N_sh0_0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   n2, n3, n5, n6, n1, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign B[31] = B[16];
  assign B[30] = B[16];
  assign B[29] = B[16];
  assign B[28] = B[16];
  assign B[27] = B[16];
  assign B[26] = B[16];
  assign B[25] = B[16];
  assign B[24] = B[16];
  assign B[23] = B[16];
  assign B[22] = B[16];
  assign B[21] = B[16];
  assign B[20] = B[16];
  assign B[19] = B[16];
  assign B[18] = B[16];
  assign B[17] = B[16];

  XOR2_X1 U26 ( .A(sel[1]), .B(sel[0]), .Z(n6) );
  CLKBUF_X3 U3 ( .A(n7), .Z(B[16]) );
  XNOR2_X2 U4 ( .A(n59), .B(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(n59), .ZN(n60) );
  BUF_X1 U6 ( .A(n62), .Z(n58) );
  XNOR2_X1 U7 ( .A(n61), .B(n58), .ZN(n1) );
  BUF_X1 U8 ( .A(n62), .Z(n57) );
  NOR2_X1 U9 ( .A1(n27), .A2(n9), .ZN(n47) );
  NOR2_X1 U10 ( .A1(n29), .A2(n9), .ZN(n48) );
  NOR2_X1 U11 ( .A1(n19), .A2(n9), .ZN(n43) );
  NOR2_X1 U12 ( .A1(n35), .A2(n9), .ZN(n51) );
  NOR2_X1 U13 ( .A1(n13), .A2(n9), .ZN(n40) );
  NOR2_X1 U14 ( .A1(n21), .A2(n9), .ZN(n44) );
  NOR2_X1 U15 ( .A1(n9), .A2(n10), .ZN(n39) );
  NOR2_X1 U16 ( .A1(n37), .A2(n9), .ZN(n52) );
  NOR2_X1 U17 ( .A1(n25), .A2(n9), .ZN(n46) );
  NOR2_X1 U18 ( .A1(n17), .A2(n9), .ZN(n42) );
  NOR2_X1 U19 ( .A1(n33), .A2(n9), .ZN(n50) );
  NOR2_X1 U20 ( .A1(n31), .A2(n9), .ZN(n49) );
  NOR2_X1 U21 ( .A1(n15), .A2(n9), .ZN(n41) );
  NOR2_X1 U22 ( .A1(n23), .A2(n9), .ZN(n45) );
  NOR2_X1 U23 ( .A1(n38), .A2(n9), .ZN(n53) );
  INV_X1 U24 ( .A(n2), .ZN(B[0]) );
  AOI22_X1 U25 ( .A1(n3), .A2(AS), .B1(n63), .B2(n5), .ZN(n2) );
  INV_X1 U27 ( .A(n3), .ZN(n5) );
  NAND2_X1 U28 ( .A1(n6), .A2(A[0]), .ZN(n3) );
  OAI21_X1 U29 ( .B1(n58), .B2(n61), .A(sel[0]), .ZN(n54) );
  INV_X1 U30 ( .A(n56), .ZN(n7) );
  NAND2_X1 U31 ( .A1(n1), .A2(n54), .ZN(n55) );
  AOI22_X1 U32 ( .A1(n58), .A2(n61), .B1(sel[0]), .B2(n1), .ZN(n8) );
  XOR2_X1 U33 ( .A(n59), .B(n64), .Z(n10) );
  XOR2_X1 U34 ( .A(n58), .B(A[1]), .Z(n11) );
  XOR2_X1 U35 ( .A(n57), .B(A[2]), .Z(n12) );
  XOR2_X1 U36 ( .A(n60), .B(A[1]), .Z(n13) );
  XOR2_X1 U37 ( .A(n57), .B(A[3]), .Z(n14) );
  XOR2_X1 U38 ( .A(n60), .B(A[2]), .Z(n15) );
  XOR2_X1 U39 ( .A(n57), .B(A[4]), .Z(n16) );
  XOR2_X1 U40 ( .A(n60), .B(A[3]), .Z(n17) );
  XOR2_X1 U41 ( .A(n58), .B(A[5]), .Z(n18) );
  XOR2_X1 U42 ( .A(n60), .B(A[4]), .Z(n19) );
  XOR2_X1 U43 ( .A(n58), .B(A[6]), .Z(n20) );
  XOR2_X1 U44 ( .A(n60), .B(A[5]), .Z(n21) );
  XOR2_X1 U45 ( .A(n58), .B(A[7]), .Z(n22) );
  XOR2_X1 U46 ( .A(n60), .B(A[6]), .Z(n23) );
  XOR2_X1 U47 ( .A(n58), .B(A[8]), .Z(n24) );
  XOR2_X1 U48 ( .A(n60), .B(A[7]), .Z(n25) );
  XOR2_X1 U49 ( .A(n58), .B(A[9]), .Z(n26) );
  XOR2_X1 U50 ( .A(n60), .B(A[8]), .Z(n27) );
  XOR2_X1 U51 ( .A(n58), .B(A[10]), .Z(n28) );
  XOR2_X1 U52 ( .A(n60), .B(A[9]), .Z(n29) );
  XOR2_X1 U53 ( .A(n58), .B(A[11]), .Z(n30) );
  XOR2_X1 U54 ( .A(n60), .B(A[10]), .Z(n31) );
  XOR2_X1 U55 ( .A(n58), .B(A[12]), .Z(n32) );
  XOR2_X1 U56 ( .A(n60), .B(A[11]), .Z(n33) );
  XOR2_X1 U57 ( .A(n58), .B(A[13]), .Z(n34) );
  XOR2_X1 U58 ( .A(n60), .B(A[12]), .Z(n35) );
  XOR2_X1 U59 ( .A(n58), .B(A[14]), .Z(n36) );
  XOR2_X1 U60 ( .A(sel[1]), .B(A[13]), .Z(n37) );
  XOR2_X1 U61 ( .A(sel[1]), .B(A[14]), .Z(n38) );
  MUX2_X1 U62 ( .A(n39), .B(n11), .S(n4), .Z(B[1]) );
  MUX2_X1 U63 ( .A(n40), .B(n12), .S(n4), .Z(B[2]) );
  MUX2_X1 U64 ( .A(n41), .B(n14), .S(n4), .Z(B[3]) );
  MUX2_X1 U65 ( .A(n42), .B(n16), .S(n4), .Z(B[4]) );
  MUX2_X1 U66 ( .A(n43), .B(n18), .S(n4), .Z(B[5]) );
  MUX2_X1 U67 ( .A(n44), .B(n20), .S(n4), .Z(B[6]) );
  MUX2_X1 U68 ( .A(n45), .B(n22), .S(n4), .Z(B[7]) );
  MUX2_X1 U69 ( .A(n46), .B(n24), .S(n4), .Z(B[8]) );
  MUX2_X1 U70 ( .A(n47), .B(n26), .S(n4), .Z(B[9]) );
  MUX2_X1 U71 ( .A(n48), .B(n28), .S(n4), .Z(B[10]) );
  MUX2_X1 U72 ( .A(n49), .B(n30), .S(n4), .Z(B[11]) );
  MUX2_X1 U73 ( .A(n50), .B(n32), .S(n4), .Z(B[12]) );
  MUX2_X1 U74 ( .A(n51), .B(n34), .S(n4), .Z(B[13]) );
  MUX2_X1 U75 ( .A(n52), .B(n36), .S(n4), .Z(B[14]) );
  MUX2_X1 U76 ( .A(n53), .B(n1), .S(n4), .Z(B[15]) );
  MUX2_X1 U77 ( .A(n8), .B(n55), .S(sel[1]), .Z(n56) );
  INV_X1 U78 ( .A(sel[1]), .ZN(n59) );
  XOR2_X2 U79 ( .A(n59), .B(n58), .Z(n9) );
  INV_X1 U80 ( .A(A[15]), .ZN(n61) );
  AOI21_X1 U81 ( .B1(sel[1]), .B2(sel[0]), .A(n63), .ZN(AS) );
  INV_X1 U82 ( .A(sel[2]), .ZN(n63) );
  INV_X1 U83 ( .A(n63), .ZN(n62) );
  INV_X1 U84 ( .A(A[0]), .ZN(n64) );
endmodule


module sum_gen_Nrca4_NB32_8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_71 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_70 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_69 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_68 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_67 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_66 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_65 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_64 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_8 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   n9, n10, g0temp, \matrixProp[0][31] , \matrixProp[0][30] ,
         \matrixProp[0][29] , \matrixProp[0][28] , \matrixProp[0][27] ,
         \matrixProp[0][26] , \matrixProp[0][25] , \matrixProp[0][24] ,
         \matrixProp[0][23] , \matrixProp[0][22] , \matrixProp[0][21] ,
         \matrixProp[0][20] , \matrixProp[0][19] , \matrixProp[0][18] ,
         \matrixProp[0][17] , \matrixProp[0][16] , \matrixProp[0][15] ,
         \matrixProp[0][14] , \matrixProp[0][13] , \matrixProp[0][12] ,
         \matrixProp[0][11] , \matrixProp[0][10] , \matrixProp[0][9] ,
         \matrixProp[0][8] , \matrixProp[0][7] , \matrixProp[0][6] ,
         \matrixProp[0][5] , \matrixProp[0][4] , \matrixProp[0][3] ,
         \matrixProp[0][2] , \matrixProp[0][1] , \matrixProp[0][0] ,
         \matrixProp[1][31] , \matrixProp[1][29] , \matrixProp[1][27] ,
         \matrixProp[1][25] , \matrixProp[1][23] , \matrixProp[1][21] ,
         \matrixProp[1][19] , \matrixProp[1][17] , \matrixProp[1][15] ,
         \matrixProp[1][13] , \matrixProp[1][11] , \matrixProp[1][9] ,
         \matrixProp[1][7] , \matrixProp[1][5] , \matrixProp[1][3] ,
         \matrixProp[2][31] , \matrixProp[2][27] , \matrixProp[2][23] ,
         \matrixProp[2][19] , \matrixProp[2][15] , \matrixProp[2][11] ,
         \matrixProp[2][7] , \matrixProp[3][31] , \matrixProp[3][23] ,
         \matrixProp[3][15] , \matrixProp[4][31] , \matrixProp[4][27] ,
         \matrixGen[0][31] , \matrixGen[0][30] , \matrixGen[0][29] ,
         \matrixGen[0][28] , \matrixGen[0][27] , \matrixGen[0][26] ,
         \matrixGen[0][25] , \matrixGen[0][24] , \matrixGen[0][23] ,
         \matrixGen[0][22] , \matrixGen[0][21] , \matrixGen[0][20] ,
         \matrixGen[0][19] , \matrixGen[0][18] , \matrixGen[0][17] ,
         \matrixGen[0][16] , \matrixGen[0][15] , \matrixGen[0][14] ,
         \matrixGen[0][13] , \matrixGen[0][12] , \matrixGen[0][11] ,
         \matrixGen[0][10] , \matrixGen[0][9] , \matrixGen[0][8] ,
         \matrixGen[0][7] , \matrixGen[0][6] , \matrixGen[0][5] ,
         \matrixGen[0][4] , \matrixGen[0][3] , \matrixGen[0][2] ,
         \matrixGen[0][1] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n1, n2, n5, n7, n8, n6;

  CLKBUF_X1 U2 ( .A(C[3]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n10), .Z(C[0]) );
  CLKBUF_X1 U4 ( .A(n1), .Z(C[1]) );
  CLKBUF_X1 U5 ( .A(\matrixGen[2][11] ), .Z(n5) );
  INV_X1 U6 ( .A(g0temp), .ZN(n7) );
  pg_net_287 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_286 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_285 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_284 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_283 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_282 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_281 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_280 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_279 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_278 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_277 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_276 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_275 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_274 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_273 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_272 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_271 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_270 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_269 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_268 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_267 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_266 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_265 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_264 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_263 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_262 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_261 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_260 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_259 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_258 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_257 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_256 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_242 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_80 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(n8), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_241 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_240 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_239 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_238 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_237 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_236 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_235 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_234 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_233 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_232 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_231 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_230 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_229 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_228 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_79 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(n10) );
  blockPG_227 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_226 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_225 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_224 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_223 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_222 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_221 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_78 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(n10), .Pik(
        \matrixProp[2][7] ), .Gij(n9) );
  blockPG_220 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_219 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_218 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_77 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(n9), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_76 gen2_4_16_2 ( .Gik(n5), .Gk_1j(n1), .Pik(\matrixProp[2][11] ), .Gij(
        C[2]) );
  blockPG_217 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_216 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_75 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(n2), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_74 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_73 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_72 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  NAND2_X1 U8 ( .A1(n6), .A2(n7), .ZN(n8) );
  NAND2_X1 U7 ( .A1(\matrixProp[0][0] ), .A2(Ci), .ZN(n6) );
  BUF_X1 U1 ( .A(n9), .Z(n1) );
endmodule


module BP_NB32_BP_LEN4_0_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  NOR4_X1 U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(EQ) );
  NAND4_X1 U2 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B[3]), .B(A[3]), .ZN(n8) );
  XNOR2_X1 U4 ( .A(B[4]), .B(A[4]), .ZN(n7) );
  XNOR2_X1 U5 ( .A(B[5]), .B(A[5]), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B[6]), .B(A[6]), .ZN(n5) );
  NAND4_X1 U7 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  OAI22_X1 U8 ( .A1(n13), .A2(n14), .B1(B[1]), .B2(n13), .ZN(n12) );
  INV_X1 U9 ( .A(A[1]), .ZN(n14) );
  AND2_X1 U10 ( .A1(B[0]), .A2(n15), .ZN(n13) );
  OAI22_X1 U11 ( .A1(A[1]), .A2(n16), .B1(n16), .B2(n17), .ZN(n11) );
  INV_X1 U12 ( .A(B[1]), .ZN(n17) );
  NOR2_X1 U13 ( .A1(n15), .A2(B[0]), .ZN(n16) );
  INV_X1 U14 ( .A(A[0]), .ZN(n15) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n10) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n2) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n1) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule


module BP_NB32_BP_LEN4_0_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n28, n30, n31, n9, n8, n7, n6, n5, n4, n34, n33, n32, n3, n29, n27,
         n26, n25, n24, n23, n22, n21, n20, n2, net413673, net413672, n50, n48,
         n47, n42, n40, n39, n19, n18, n17, n16, n15, n1, n41, n14, n13, n12,
         n11, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60;

  AND2_X1 U31 ( .A1(B[0]), .A2(n30), .ZN(n28) );
  NOR2_X1 U34 ( .A1(n30), .A2(B[0]), .ZN(n31) );
  INV_X1 U35 ( .A(A[0]), .ZN(n30) );
  XNOR2_X1 U5 ( .A(B[11]), .B(A[11]), .ZN(n2) );
  XNOR2_X1 U6 ( .A(B[12]), .B(A[12]), .ZN(n3) );
  XNOR2_X1 U7 ( .A(B[13]), .B(A[13]), .ZN(n4) );
  XNOR2_X1 U8 ( .A(B[14]), .B(A[14]), .ZN(n5) );
  AND4_X1 U4 ( .A1(n2), .A2(n3), .A3(n4), .A4(n5), .ZN(n33) );
  AND2_X1 U10 ( .A1(n33), .A2(n34), .ZN(n7) );
  XNOR2_X1 U37 ( .A(B[2]), .B(A[2]), .ZN(n24) );
  XNOR2_X1 U36 ( .A(B[31]), .B(A[31]), .ZN(n25) );
  INV_X1 U33 ( .A(B[1]), .ZN(n32) );
  OAI22_X1 U32 ( .A1(A[1]), .A2(n31), .B1(n31), .B2(n32), .ZN(n26) );
  INV_X1 U30 ( .A(A[1]), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n28), .A2(n29), .B1(B[1]), .B2(n28), .ZN(n27) );
  AND4_X1 U11 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n8) );
  XNOR2_X1 U28 ( .A(B[6]), .B(A[6]), .ZN(n20) );
  XNOR2_X1 U27 ( .A(B[5]), .B(A[5]), .ZN(n21) );
  XNOR2_X1 U26 ( .A(B[4]), .B(A[4]), .ZN(n22) );
  XNOR2_X1 U25 ( .A(B[3]), .B(A[3]), .ZN(n23) );
  AND4_X1 U12 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n9) );
  NAND3_X1 U9 ( .A1(n7), .A2(n8), .A3(n9), .ZN(n6) );
  XNOR2_X1 U23 ( .A(B[29]), .B(A[29]), .ZN(n17) );
  XNOR2_X1 U24 ( .A(B[30]), .B(A[30]), .ZN(n18) );
  XNOR2_X1 U21 ( .A(B[27]), .B(A[27]), .ZN(n15) );
  XNOR2_X1 U22 ( .A(B[28]), .B(A[28]), .ZN(n16) );
  AND4_X1 U20 ( .A1(n17), .A2(n18), .A3(n15), .A4(n16), .ZN(n39) );
  XOR2_X1 U50 ( .A(B[24]), .B(A[24]), .Z(n48) );
  INV_X2 syn33 ( .A(n48), .ZN(net413673) );
  INV_X1 U2 ( .A(A[26]), .ZN(n1) );
  XNOR2_X1 U3 ( .A(B[26]), .B(n1), .ZN(n50) );
  NOR2_X1 U19 ( .A1(n19), .A2(n6), .ZN(EQ) );
  XNOR2_X1 U17 ( .A(B[21]), .B(A[21]), .ZN(n13) );
  XNOR2_X1 U18 ( .A(B[22]), .B(A[22]), .ZN(n14) );
  XNOR2_X1 U15 ( .A(B[19]), .B(A[19]), .ZN(n11) );
  XNOR2_X1 U16 ( .A(B[20]), .B(A[20]), .ZN(n12) );
  NAND4_X1 U43 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(n19) );
  AND4_X1 U14 ( .A1(n13), .A2(n14), .A3(n11), .A4(n12), .ZN(n41) );
  AND4_X1 U1 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(n34) );
  XNOR2_X1 U13 ( .A(B[7]), .B(A[7]), .ZN(n51) );
  XNOR2_X1 U38 ( .A(B[8]), .B(A[8]), .ZN(n52) );
  XNOR2_X1 U39 ( .A(B[9]), .B(A[9]), .ZN(n53) );
  XNOR2_X1 U40 ( .A(B[10]), .B(A[10]), .ZN(n54) );
  AND4_X1 U41 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(n42) );
  XNOR2_X1 U42 ( .A(B[15]), .B(A[15]), .ZN(n55) );
  XNOR2_X1 U44 ( .A(B[16]), .B(A[16]), .ZN(n56) );
  XNOR2_X1 U45 ( .A(B[17]), .B(A[17]), .ZN(n57) );
  XNOR2_X1 U46 ( .A(B[18]), .B(A[18]), .ZN(n58) );
  AND3_X1 U47 ( .A1(net413672), .A2(n59), .A3(net413673), .ZN(n40) );
  NOR2_X1 U48 ( .A1(n50), .A2(n47), .ZN(n59) );
  XNOR2_X1 U49 ( .A(B[23]), .B(n60), .ZN(n47) );
  INV_X32 U51 ( .A(A[23]), .ZN(n60) );
  XNOR2_X1 U52 ( .A(B[25]), .B(A[25]), .ZN(net413672) );
endmodule


module FD_NB5_0 ( CK, RESET, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
endmodule


module EXECUTION_UNIT_NB32_LS5_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , n1;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XNOR2_X1 U1 ( .A(A[31]), .B(n1), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n1) );
  XOR2_X1 U3 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  AND2_X1 U4 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  XOR2_X1 U5 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  AND2_X1 U6 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  XOR2_X1 U7 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  AND2_X1 U8 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  XOR2_X1 U9 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  AND2_X1 U10 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  XOR2_X1 U11 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  AND2_X1 U12 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  XOR2_X1 U13 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  AND2_X1 U14 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  XOR2_X1 U15 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  AND2_X1 U16 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  XOR2_X1 U17 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  AND2_X1 U18 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  XOR2_X1 U19 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  AND2_X1 U20 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  XOR2_X1 U21 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  AND2_X1 U22 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  XOR2_X1 U23 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  AND2_X1 U24 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  XOR2_X1 U25 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  AND2_X1 U26 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  XOR2_X1 U27 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  AND2_X1 U28 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  XOR2_X1 U29 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  AND2_X1 U30 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  XOR2_X1 U31 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  AND2_X1 U32 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  XOR2_X1 U33 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  AND2_X1 U34 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  XOR2_X1 U35 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  AND2_X1 U36 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  XOR2_X1 U37 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  AND2_X1 U38 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  XOR2_X1 U39 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  AND2_X1 U40 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  XOR2_X1 U41 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  AND2_X1 U42 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  XOR2_X1 U43 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  AND2_X1 U44 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  XOR2_X1 U45 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  AND2_X1 U46 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  XOR2_X1 U47 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  AND2_X1 U48 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  XOR2_X1 U49 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  AND2_X1 U50 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  XOR2_X1 U51 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  AND2_X1 U52 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  XOR2_X1 U53 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  AND2_X1 U54 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  XOR2_X1 U55 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  AND2_X1 U56 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  XOR2_X1 U57 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  INV_X1 U58 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module MUX61_generic_NB32_0 ( A, B, C, D, E, F, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [2:0] SEL;
  output [31:0] Y;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, n2, n3, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n1, n4, n11, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95;

  DLH_X1 \Y_reg[31]  ( .G(n93), .D(N44), .Q(Y[31]) );
  DLH_X1 \Y_reg[30]  ( .G(n93), .D(N42), .Q(Y[30]) );
  DLH_X1 \Y_reg[29]  ( .G(n93), .D(N41), .Q(Y[29]) );
  DLH_X1 \Y_reg[28]  ( .G(n93), .D(N40), .Q(Y[28]) );
  DLH_X1 \Y_reg[27]  ( .G(n93), .D(N39), .Q(Y[27]) );
  DLH_X1 \Y_reg[26]  ( .G(n93), .D(N38), .Q(Y[26]) );
  DLH_X1 \Y_reg[25]  ( .G(n93), .D(N37), .Q(Y[25]) );
  DLH_X1 \Y_reg[24]  ( .G(n93), .D(N36), .Q(Y[24]) );
  DLH_X1 \Y_reg[23]  ( .G(n93), .D(N35), .Q(Y[23]) );
  DLH_X1 \Y_reg[22]  ( .G(n93), .D(N34), .Q(Y[22]) );
  DLH_X1 \Y_reg[21]  ( .G(n93), .D(N33), .Q(Y[21]) );
  DLH_X1 \Y_reg[20]  ( .G(n94), .D(N32), .Q(Y[20]) );
  DLH_X1 \Y_reg[19]  ( .G(n94), .D(N31), .Q(Y[19]) );
  DLH_X1 \Y_reg[18]  ( .G(n94), .D(N30), .Q(Y[18]) );
  DLH_X1 \Y_reg[17]  ( .G(n94), .D(N29), .Q(Y[17]) );
  DLH_X1 \Y_reg[16]  ( .G(n94), .D(N28), .Q(Y[16]) );
  DLH_X1 \Y_reg[15]  ( .G(n94), .D(N27), .Q(Y[15]) );
  DLH_X1 \Y_reg[14]  ( .G(n94), .D(N26), .Q(Y[14]) );
  DLH_X1 \Y_reg[13]  ( .G(n94), .D(N25), .Q(Y[13]) );
  DLH_X1 \Y_reg[12]  ( .G(n94), .D(N24), .Q(Y[12]) );
  DLH_X1 \Y_reg[11]  ( .G(n94), .D(N23), .Q(Y[11]) );
  DLH_X1 \Y_reg[10]  ( .G(n94), .D(N22), .Q(Y[10]) );
  DLH_X1 \Y_reg[9]  ( .G(n95), .D(N21), .Q(Y[9]) );
  DLH_X1 \Y_reg[8]  ( .G(n95), .D(N20), .Q(Y[8]) );
  DLH_X1 \Y_reg[7]  ( .G(n95), .D(N19), .Q(Y[7]) );
  DLH_X1 \Y_reg[6]  ( .G(n95), .D(N18), .Q(Y[6]) );
  DLH_X1 \Y_reg[5]  ( .G(n95), .D(N17), .Q(Y[5]) );
  DLH_X1 \Y_reg[4]  ( .G(n95), .D(N16), .Q(Y[4]) );
  DLH_X1 \Y_reg[3]  ( .G(n95), .D(N15), .Q(Y[3]) );
  DLH_X1 \Y_reg[2]  ( .G(n95), .D(N14), .Q(Y[2]) );
  DLH_X1 \Y_reg[1]  ( .G(n95), .D(N13), .Q(Y[1]) );
  DLH_X1 \Y_reg[0]  ( .G(n95), .D(N12), .Q(Y[0]) );
  NAND3_X1 U109 ( .A1(n76), .A2(n77), .A3(SEL[2]), .ZN(n10) );
  NAND3_X1 U110 ( .A1(SEL[0]), .A2(n77), .A3(SEL[2]), .ZN(n12) );
  AOI222_X4 U2 ( .A1(A[26]), .A2(n82), .B1(C[26]), .B2(n79), .C1(B[26]), .C2(
        n4), .ZN(n22) );
  BUF_X1 U3 ( .A(n5), .Z(n88) );
  BUF_X1 U4 ( .A(n5), .Z(n89) );
  BUF_X1 U5 ( .A(n6), .Z(n85) );
  BUF_X1 U6 ( .A(n6), .Z(n86) );
  BUF_X1 U7 ( .A(n5), .Z(n90) );
  BUF_X1 U8 ( .A(n6), .Z(n87) );
  BUF_X1 U9 ( .A(N43), .Z(n94) );
  BUF_X1 U10 ( .A(N43), .Z(n93) );
  BUF_X1 U11 ( .A(N43), .Z(n95) );
  INV_X1 U12 ( .A(n1), .ZN(n91) );
  INV_X1 U13 ( .A(n1), .ZN(n92) );
  BUF_X1 U14 ( .A(n7), .Z(n83) );
  BUF_X1 U15 ( .A(n8), .Z(n81) );
  BUF_X1 U16 ( .A(n9), .Z(n78) );
  BUF_X1 U17 ( .A(n8), .Z(n80) );
  BUF_X1 U18 ( .A(n9), .Z(n11) );
  BUF_X1 U19 ( .A(n7), .Z(n82) );
  BUF_X1 U20 ( .A(n8), .Z(n79) );
  BUF_X1 U21 ( .A(n9), .Z(n4) );
  BUF_X1 U22 ( .A(n7), .Z(n84) );
  NAND4_X1 U23 ( .A1(n10), .A2(n1), .A3(n12), .A4(n13), .ZN(N43) );
  NOR3_X1 U24 ( .A1(n81), .A2(n82), .A3(n4), .ZN(n13) );
  INV_X1 U25 ( .A(n12), .ZN(n5) );
  INV_X1 U26 ( .A(n10), .ZN(n6) );
  NOR3_X1 U27 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n7) );
  NOR3_X1 U28 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n77), .ZN(n8) );
  NOR3_X1 U29 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n76), .ZN(n9) );
  OR3_X1 U30 ( .A1(n76), .A2(SEL[2]), .A3(n77), .ZN(n1) );
  INV_X1 U31 ( .A(SEL[1]), .ZN(n77) );
  INV_X1 U32 ( .A(SEL[0]), .ZN(n76) );
  NAND2_X1 U33 ( .A1(n14), .A2(n15), .ZN(N42) );
  AOI222_X1 U34 ( .A1(D[30]), .A2(n91), .B1(F[30]), .B2(n90), .C1(E[30]), .C2(
        n87), .ZN(n15) );
  NAND2_X1 U35 ( .A1(n72), .A2(n73), .ZN(N13) );
  AOI222_X1 U36 ( .A1(A[1]), .A2(n84), .B1(C[1]), .B2(n81), .C1(B[1]), .C2(n78), .ZN(n72) );
  AOI222_X1 U37 ( .A1(D[1]), .A2(n91), .B1(F[1]), .B2(n88), .C1(E[1]), .C2(n85), .ZN(n73) );
  NAND2_X1 U38 ( .A1(n70), .A2(n71), .ZN(N14) );
  AOI222_X1 U39 ( .A1(A[2]), .A2(n84), .B1(C[2]), .B2(n81), .C1(B[2]), .C2(n78), .ZN(n70) );
  AOI222_X1 U40 ( .A1(D[2]), .A2(n91), .B1(F[2]), .B2(n88), .C1(E[2]), .C2(n85), .ZN(n71) );
  NAND2_X1 U41 ( .A1(n68), .A2(n69), .ZN(N15) );
  AOI222_X1 U42 ( .A1(A[3]), .A2(n84), .B1(C[3]), .B2(n81), .C1(B[3]), .C2(n78), .ZN(n68) );
  AOI222_X1 U43 ( .A1(D[3]), .A2(n91), .B1(F[3]), .B2(n88), .C1(E[3]), .C2(n85), .ZN(n69) );
  NAND2_X1 U44 ( .A1(n66), .A2(n67), .ZN(N16) );
  AOI222_X1 U45 ( .A1(A[4]), .A2(n84), .B1(C[4]), .B2(n81), .C1(B[4]), .C2(n78), .ZN(n66) );
  AOI222_X1 U46 ( .A1(D[4]), .A2(n91), .B1(F[4]), .B2(n88), .C1(E[4]), .C2(n85), .ZN(n67) );
  NAND2_X1 U47 ( .A1(n64), .A2(n65), .ZN(N17) );
  AOI222_X1 U48 ( .A1(A[5]), .A2(n84), .B1(C[5]), .B2(n81), .C1(B[5]), .C2(n78), .ZN(n64) );
  AOI222_X1 U49 ( .A1(D[5]), .A2(n91), .B1(F[5]), .B2(n88), .C1(E[5]), .C2(n85), .ZN(n65) );
  NAND2_X1 U50 ( .A1(n62), .A2(n63), .ZN(N18) );
  AOI222_X1 U51 ( .A1(A[6]), .A2(n84), .B1(C[6]), .B2(n81), .C1(B[6]), .C2(n78), .ZN(n62) );
  AOI222_X1 U52 ( .A1(D[6]), .A2(n91), .B1(F[6]), .B2(n88), .C1(E[6]), .C2(n85), .ZN(n63) );
  NAND2_X1 U53 ( .A1(n60), .A2(n61), .ZN(N19) );
  AOI222_X1 U54 ( .A1(A[7]), .A2(n84), .B1(C[7]), .B2(n81), .C1(B[7]), .C2(n78), .ZN(n60) );
  AOI222_X1 U55 ( .A1(D[7]), .A2(n91), .B1(F[7]), .B2(n88), .C1(E[7]), .C2(n85), .ZN(n61) );
  NAND2_X1 U56 ( .A1(n58), .A2(n59), .ZN(N20) );
  AOI222_X1 U57 ( .A1(A[8]), .A2(n83), .B1(C[8]), .B2(n81), .C1(B[8]), .C2(n78), .ZN(n58) );
  AOI222_X1 U58 ( .A1(D[8]), .A2(n91), .B1(F[8]), .B2(n88), .C1(E[8]), .C2(n85), .ZN(n59) );
  NAND2_X1 U59 ( .A1(n56), .A2(n57), .ZN(N21) );
  AOI222_X1 U60 ( .A1(A[9]), .A2(n83), .B1(C[9]), .B2(n80), .C1(B[9]), .C2(n78), .ZN(n56) );
  AOI222_X1 U61 ( .A1(D[9]), .A2(n91), .B1(F[9]), .B2(n88), .C1(E[9]), .C2(n85), .ZN(n57) );
  NAND2_X1 U62 ( .A1(n74), .A2(n75), .ZN(N12) );
  AOI222_X1 U63 ( .A1(A[0]), .A2(n82), .B1(C[0]), .B2(n79), .C1(B[0]), .C2(n4), 
        .ZN(n74) );
  AOI222_X1 U64 ( .A1(D[0]), .A2(n91), .B1(F[0]), .B2(n88), .C1(E[0]), .C2(n85), .ZN(n75) );
  NAND2_X1 U65 ( .A1(n54), .A2(n55), .ZN(N22) );
  AOI222_X1 U66 ( .A1(A[10]), .A2(n83), .B1(C[10]), .B2(n80), .C1(B[10]), .C2(
        n11), .ZN(n54) );
  AOI222_X1 U67 ( .A1(D[10]), .A2(n91), .B1(F[10]), .B2(n88), .C1(E[10]), .C2(
        n85), .ZN(n55) );
  NAND2_X1 U68 ( .A1(n52), .A2(n53), .ZN(N23) );
  AOI222_X1 U69 ( .A1(A[11]), .A2(n83), .B1(C[11]), .B2(n80), .C1(B[11]), .C2(
        n11), .ZN(n52) );
  AOI222_X1 U70 ( .A1(D[11]), .A2(n91), .B1(F[11]), .B2(n88), .C1(E[11]), .C2(
        n85), .ZN(n53) );
  NAND2_X1 U71 ( .A1(n50), .A2(n51), .ZN(N24) );
  AOI222_X1 U72 ( .A1(A[12]), .A2(n83), .B1(C[12]), .B2(n80), .C1(B[12]), .C2(
        n11), .ZN(n50) );
  AOI222_X1 U73 ( .A1(D[12]), .A2(n92), .B1(F[12]), .B2(n89), .C1(E[12]), .C2(
        n86), .ZN(n51) );
  NAND2_X1 U74 ( .A1(n48), .A2(n49), .ZN(N25) );
  AOI222_X1 U75 ( .A1(A[13]), .A2(n83), .B1(C[13]), .B2(n80), .C1(B[13]), .C2(
        n11), .ZN(n48) );
  AOI222_X1 U76 ( .A1(D[13]), .A2(n92), .B1(F[13]), .B2(n89), .C1(E[13]), .C2(
        n86), .ZN(n49) );
  NAND2_X1 U77 ( .A1(n46), .A2(n47), .ZN(N26) );
  AOI222_X1 U78 ( .A1(A[14]), .A2(n83), .B1(C[14]), .B2(n80), .C1(B[14]), .C2(
        n11), .ZN(n46) );
  AOI222_X1 U79 ( .A1(D[14]), .A2(n92), .B1(F[14]), .B2(n89), .C1(E[14]), .C2(
        n86), .ZN(n47) );
  NAND2_X1 U80 ( .A1(n44), .A2(n45), .ZN(N27) );
  AOI222_X1 U81 ( .A1(A[15]), .A2(n83), .B1(C[15]), .B2(n80), .C1(B[15]), .C2(
        n11), .ZN(n44) );
  AOI222_X1 U82 ( .A1(D[15]), .A2(n92), .B1(F[15]), .B2(n89), .C1(E[15]), .C2(
        n86), .ZN(n45) );
  NAND2_X1 U83 ( .A1(n42), .A2(n43), .ZN(N28) );
  AOI222_X1 U84 ( .A1(A[16]), .A2(n83), .B1(C[16]), .B2(n80), .C1(B[16]), .C2(
        n11), .ZN(n42) );
  AOI222_X1 U85 ( .A1(D[16]), .A2(n92), .B1(F[16]), .B2(n89), .C1(E[16]), .C2(
        n86), .ZN(n43) );
  NAND2_X1 U86 ( .A1(n40), .A2(n41), .ZN(N29) );
  AOI222_X1 U87 ( .A1(A[17]), .A2(n83), .B1(C[17]), .B2(n80), .C1(B[17]), .C2(
        n11), .ZN(n40) );
  AOI222_X1 U88 ( .A1(D[17]), .A2(n92), .B1(F[17]), .B2(n89), .C1(E[17]), .C2(
        n86), .ZN(n41) );
  NAND2_X1 U89 ( .A1(n38), .A2(n39), .ZN(N30) );
  AOI222_X1 U90 ( .A1(A[18]), .A2(n83), .B1(C[18]), .B2(n80), .C1(B[18]), .C2(
        n11), .ZN(n38) );
  AOI222_X1 U91 ( .A1(D[18]), .A2(n92), .B1(F[18]), .B2(n89), .C1(E[18]), .C2(
        n86), .ZN(n39) );
  NAND2_X1 U92 ( .A1(n36), .A2(n37), .ZN(N31) );
  AOI222_X1 U93 ( .A1(A[19]), .A2(n83), .B1(C[19]), .B2(n80), .C1(B[19]), .C2(
        n11), .ZN(n36) );
  AOI222_X1 U94 ( .A1(D[19]), .A2(n92), .B1(F[19]), .B2(n89), .C1(E[19]), .C2(
        n86), .ZN(n37) );
  NAND2_X1 U95 ( .A1(n34), .A2(n35), .ZN(N32) );
  AOI222_X1 U96 ( .A1(A[20]), .A2(n82), .B1(C[20]), .B2(n79), .C1(B[20]), .C2(
        n11), .ZN(n34) );
  AOI222_X1 U97 ( .A1(D[20]), .A2(n92), .B1(F[20]), .B2(n89), .C1(E[20]), .C2(
        n86), .ZN(n35) );
  NAND2_X1 U98 ( .A1(n30), .A2(n31), .ZN(N34) );
  AOI222_X1 U100 ( .A1(D[22]), .A2(n92), .B1(F[22]), .B2(n89), .C1(E[22]), 
        .C2(n86), .ZN(n31) );
  NAND2_X1 U101 ( .A1(n28), .A2(n29), .ZN(N35) );
  AOI222_X1 U102 ( .A1(A[23]), .A2(n82), .B1(C[23]), .B2(n79), .C1(B[23]), 
        .C2(n4), .ZN(n28) );
  AOI222_X1 U103 ( .A1(D[23]), .A2(n92), .B1(F[23]), .B2(n89), .C1(E[23]), 
        .C2(n86), .ZN(n29) );
  NAND2_X1 U104 ( .A1(n26), .A2(n27), .ZN(N36) );
  AOI222_X1 U105 ( .A1(A[24]), .A2(n82), .B1(C[24]), .B2(n79), .C1(B[24]), 
        .C2(n4), .ZN(n26) );
  AOI222_X1 U106 ( .A1(D[24]), .A2(n92), .B1(F[24]), .B2(n90), .C1(E[24]), 
        .C2(n87), .ZN(n27) );
  NAND2_X1 U107 ( .A1(n22), .A2(n23), .ZN(N38) );
  AOI222_X1 U108 ( .A1(D[26]), .A2(n91), .B1(F[26]), .B2(n90), .C1(E[26]), 
        .C2(n87), .ZN(n23) );
  NAND2_X1 U111 ( .A1(n20), .A2(n21), .ZN(N39) );
  AOI222_X1 U112 ( .A1(A[27]), .A2(n82), .B1(C[27]), .B2(n79), .C1(B[27]), 
        .C2(n4), .ZN(n20) );
  AOI222_X1 U113 ( .A1(D[27]), .A2(n92), .B1(F[27]), .B2(n90), .C1(E[27]), 
        .C2(n87), .ZN(n21) );
  NAND2_X1 U114 ( .A1(n18), .A2(n19), .ZN(N40) );
  AOI222_X1 U115 ( .A1(A[28]), .A2(n82), .B1(C[28]), .B2(n79), .C1(B[28]), 
        .C2(n4), .ZN(n18) );
  AOI222_X1 U116 ( .A1(D[28]), .A2(n91), .B1(F[28]), .B2(n90), .C1(E[28]), 
        .C2(n87), .ZN(n19) );
  NAND2_X1 U117 ( .A1(n2), .A2(n3), .ZN(N44) );
  AOI222_X1 U118 ( .A1(A[31]), .A2(n83), .B1(C[31]), .B2(n80), .C1(B[31]), 
        .C2(n11), .ZN(n2) );
  AOI222_X1 U119 ( .A1(D[31]), .A2(n92), .B1(F[31]), .B2(n90), .C1(E[31]), 
        .C2(n87), .ZN(n3) );
  NAND2_X1 U120 ( .A1(n24), .A2(n25), .ZN(N37) );
  AOI222_X1 U121 ( .A1(A[25]), .A2(n82), .B1(C[25]), .B2(n79), .C1(B[25]), 
        .C2(n4), .ZN(n24) );
  AOI222_X1 U122 ( .A1(D[25]), .A2(n91), .B1(F[25]), .B2(n90), .C1(E[25]), 
        .C2(n87), .ZN(n25) );
  NAND2_X1 U123 ( .A1(n16), .A2(n17), .ZN(N41) );
  AOI222_X1 U124 ( .A1(A[29]), .A2(n82), .B1(C[29]), .B2(n79), .C1(B[29]), 
        .C2(n4), .ZN(n16) );
  AOI222_X1 U125 ( .A1(D[29]), .A2(n92), .B1(F[29]), .B2(n90), .C1(E[29]), 
        .C2(n87), .ZN(n17) );
  NAND2_X1 U126 ( .A1(n32), .A2(n33), .ZN(N33) );
  AOI222_X1 U127 ( .A1(A[21]), .A2(n82), .B1(C[21]), .B2(n79), .C1(B[21]), 
        .C2(n4), .ZN(n32) );
  AOI222_X1 U128 ( .A1(D[21]), .A2(n92), .B1(F[21]), .B2(n89), .C1(E[21]), 
        .C2(n86), .ZN(n33) );
  AOI222_X1 U129 ( .A1(A[30]), .A2(n82), .B1(C[30]), .B2(n79), .C1(B[30]), 
        .C2(n4), .ZN(n14) );
  AOI222_X1 U99 ( .A1(A[22]), .A2(n82), .B1(C[22]), .B2(n79), .C1(B[22]), .C2(
        n4), .ZN(n30) );
endmodule


module FD_NB32_3 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n33, n34, n35;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n35), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n35), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n34), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n34), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n34), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n34), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n33), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n33), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n33), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n33), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n33), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n33), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n33), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n33), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n33), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n33), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n33), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n33), .Q(Q[0]) );
  BUF_X1 U3 ( .A(RESET), .Z(n33) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
endmodule


module FD_NB5_1 ( CK, RESET, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET;


  SDFFR_X1 \TMP_Q_reg[1]  ( .D(1'b0), .SI(D[1]), .SE(1'b1), .CK(CK), .RN(RESET), .Q(Q[1]) );
  SDFFR_X1 \TMP_Q_reg[2]  ( .D(1'b0), .SI(D[2]), .SE(1'b1), .CK(CK), .RN(RESET), .Q(Q[2]) );
  SDFFR_X1 \TMP_Q_reg[4]  ( .D(1'b0), .SI(D[4]), .SE(1'b1), .CK(CK), .RN(RESET), .Q(Q[4]) );
  SDFFR_X1 \TMP_Q_reg[3]  ( .D(1'b0), .SI(D[3]), .SE(1'b1), .CK(CK), .RN(RESET), .Q(Q[3]) );
  SDFFR_X1 \TMP_Q_reg[0]  ( .D(1'b0), .SI(D[0]), .SE(1'b1), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module LOGIC_NB32_0 ( SEL, A, B, RES );
  input [3:0] SEL;
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  wire   n65, n67, n69, n70, n71, n73, n75, n77, n78, n79, n81, n83, n85, n87,
         n89, n91, n93, n94, n95, n96, n97, n98, n99, n100, n101, n103, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n147, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n169, n170, n171, n173, n175, n177,
         n178, n179, n181, n183, n185, n186, n187, n189, n191, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38;

  INV_X1 U1 ( .A(A[31]), .ZN(n96) );
  INV_X1 U2 ( .A(A[28]), .ZN(n112) );
  INV_X1 U3 ( .A(A[25]), .ZN(n124) );
  INV_X1 U4 ( .A(A[26]), .ZN(n120) );
  INV_X1 U5 ( .A(A[29]), .ZN(n108) );
  INV_X1 U6 ( .A(A[18]), .ZN(n156) );
  INV_X1 U7 ( .A(A[21]), .ZN(n140) );
  INV_X1 U8 ( .A(A[20]), .ZN(n144) );
  INV_X1 U9 ( .A(A[24]), .ZN(n128) );
  INV_X1 U10 ( .A(A[19]), .ZN(n152) );
  INV_X1 U11 ( .A(A[27]), .ZN(n116) );
  AOI22_X1 U12 ( .A1(n27), .A2(n22), .B1(A[10]), .B2(n33), .ZN(n187) );
  AOI22_X1 U13 ( .A1(n30), .A2(n22), .B1(A[10]), .B2(n36), .ZN(n185) );
  AOI22_X1 U14 ( .A1(n27), .A2(n24), .B1(A[12]), .B2(n33), .ZN(n179) );
  AOI22_X1 U15 ( .A1(n30), .A2(n24), .B1(A[12]), .B2(n36), .ZN(n177) );
  AOI22_X1 U16 ( .A1(n28), .A2(n14), .B1(A[2]), .B2(n34), .ZN(n103) );
  AOI22_X1 U17 ( .A1(n31), .A2(n14), .B1(A[2]), .B2(n37), .ZN(n101) );
  AOI22_X1 U18 ( .A1(n27), .A2(n23), .B1(A[11]), .B2(n33), .ZN(n183) );
  AOI22_X1 U19 ( .A1(n30), .A2(n23), .B1(A[11]), .B2(n36), .ZN(n181) );
  AOI22_X1 U20 ( .A1(n27), .A2(n25), .B1(A[13]), .B2(n33), .ZN(n175) );
  AOI22_X1 U21 ( .A1(n30), .A2(n25), .B1(A[13]), .B2(n36), .ZN(n173) );
  INV_X1 U22 ( .A(A[16]), .ZN(n164) );
  INV_X1 U23 ( .A(A[23]), .ZN(n132) );
  OAI22_X1 U24 ( .A1(n93), .A2(n94), .B1(B[31]), .B2(n95), .ZN(RES[31]) );
  INV_X1 U25 ( .A(B[31]), .ZN(n94) );
  AOI22_X1 U26 ( .A1(n32), .A2(n96), .B1(A[31]), .B2(n38), .ZN(n93) );
  AOI22_X1 U27 ( .A1(n29), .A2(n96), .B1(A[31]), .B2(n35), .ZN(n95) );
  INV_X1 U28 ( .A(A[30]), .ZN(n100) );
  OAI22_X1 U29 ( .A1(n109), .A2(n110), .B1(B[28]), .B2(n111), .ZN(RES[28]) );
  INV_X1 U30 ( .A(B[28]), .ZN(n110) );
  AOI22_X1 U31 ( .A1(n31), .A2(n112), .B1(A[28]), .B2(n37), .ZN(n109) );
  AOI22_X1 U32 ( .A1(n28), .A2(n112), .B1(A[28]), .B2(n34), .ZN(n111) );
  OAI22_X1 U33 ( .A1(n121), .A2(n122), .B1(B[25]), .B2(n123), .ZN(RES[25]) );
  INV_X1 U34 ( .A(B[25]), .ZN(n122) );
  AOI22_X1 U35 ( .A1(n31), .A2(n124), .B1(A[25]), .B2(n37), .ZN(n121) );
  AOI22_X1 U36 ( .A1(n28), .A2(n124), .B1(A[25]), .B2(n34), .ZN(n123) );
  OAI22_X1 U37 ( .A1(n117), .A2(n118), .B1(B[26]), .B2(n119), .ZN(RES[26]) );
  INV_X1 U38 ( .A(B[26]), .ZN(n118) );
  AOI22_X1 U39 ( .A1(n31), .A2(n120), .B1(A[26]), .B2(n37), .ZN(n117) );
  AOI22_X1 U40 ( .A1(n28), .A2(n120), .B1(A[26]), .B2(n34), .ZN(n119) );
  OAI22_X1 U41 ( .A1(n105), .A2(n106), .B1(B[29]), .B2(n107), .ZN(RES[29]) );
  INV_X1 U42 ( .A(B[29]), .ZN(n106) );
  AOI22_X1 U43 ( .A1(n31), .A2(n108), .B1(A[29]), .B2(n37), .ZN(n105) );
  AOI22_X1 U44 ( .A1(n28), .A2(n108), .B1(A[29]), .B2(n34), .ZN(n107) );
  OAI22_X1 U45 ( .A1(n153), .A2(n154), .B1(B[18]), .B2(n155), .ZN(RES[18]) );
  INV_X1 U46 ( .A(B[18]), .ZN(n154) );
  AOI22_X1 U47 ( .A1(n30), .A2(n156), .B1(A[18]), .B2(n36), .ZN(n153) );
  AOI22_X1 U48 ( .A1(n27), .A2(n156), .B1(A[18]), .B2(n33), .ZN(n155) );
  OAI22_X1 U49 ( .A1(n137), .A2(n138), .B1(B[21]), .B2(n139), .ZN(RES[21]) );
  INV_X1 U50 ( .A(B[21]), .ZN(n138) );
  AOI22_X1 U51 ( .A1(n31), .A2(n140), .B1(A[21]), .B2(n37), .ZN(n137) );
  AOI22_X1 U52 ( .A1(n28), .A2(n140), .B1(A[21]), .B2(n34), .ZN(n139) );
  OAI22_X1 U53 ( .A1(n141), .A2(n142), .B1(B[20]), .B2(n143), .ZN(RES[20]) );
  INV_X1 U54 ( .A(B[20]), .ZN(n142) );
  AOI22_X1 U55 ( .A1(n31), .A2(n144), .B1(A[20]), .B2(n37), .ZN(n141) );
  AOI22_X1 U56 ( .A1(n28), .A2(n144), .B1(A[20]), .B2(n34), .ZN(n143) );
  OAI22_X1 U57 ( .A1(n125), .A2(n126), .B1(B[24]), .B2(n127), .ZN(RES[24]) );
  INV_X1 U58 ( .A(B[24]), .ZN(n126) );
  AOI22_X1 U59 ( .A1(n31), .A2(n128), .B1(A[24]), .B2(n37), .ZN(n125) );
  AOI22_X1 U60 ( .A1(n28), .A2(n128), .B1(A[24]), .B2(n34), .ZN(n127) );
  OAI22_X1 U61 ( .A1(n149), .A2(n150), .B1(B[19]), .B2(n151), .ZN(RES[19]) );
  INV_X1 U62 ( .A(B[19]), .ZN(n150) );
  AOI22_X1 U63 ( .A1(n30), .A2(n152), .B1(A[19]), .B2(n36), .ZN(n149) );
  AOI22_X1 U64 ( .A1(n27), .A2(n152), .B1(A[19]), .B2(n33), .ZN(n151) );
  OAI22_X1 U65 ( .A1(n113), .A2(n114), .B1(B[27]), .B2(n115), .ZN(RES[27]) );
  INV_X1 U66 ( .A(B[27]), .ZN(n114) );
  AOI22_X1 U67 ( .A1(n31), .A2(n116), .B1(A[27]), .B2(n37), .ZN(n113) );
  AOI22_X1 U68 ( .A1(n28), .A2(n116), .B1(A[27]), .B2(n34), .ZN(n115) );
  OAI22_X1 U69 ( .A1(n161), .A2(n162), .B1(B[16]), .B2(n163), .ZN(RES[16]) );
  INV_X1 U70 ( .A(B[16]), .ZN(n162) );
  AOI22_X1 U71 ( .A1(n30), .A2(n164), .B1(A[16]), .B2(n36), .ZN(n161) );
  AOI22_X1 U72 ( .A1(n27), .A2(n164), .B1(A[16]), .B2(n33), .ZN(n163) );
  OAI22_X1 U73 ( .A1(n129), .A2(n130), .B1(B[23]), .B2(n131), .ZN(RES[23]) );
  INV_X1 U74 ( .A(B[23]), .ZN(n130) );
  AOI22_X1 U75 ( .A1(n31), .A2(n132), .B1(A[23]), .B2(n37), .ZN(n129) );
  AOI22_X1 U76 ( .A1(n28), .A2(n132), .B1(A[23]), .B2(n34), .ZN(n131) );
  OAI22_X1 U77 ( .A1(n157), .A2(n158), .B1(B[17]), .B2(n159), .ZN(RES[17]) );
  INV_X1 U78 ( .A(B[17]), .ZN(n158) );
  OAI22_X1 U79 ( .A1(n133), .A2(n134), .B1(B[22]), .B2(n135), .ZN(RES[22]) );
  INV_X1 U80 ( .A(B[22]), .ZN(n134) );
  OAI22_X1 U81 ( .A1(n97), .A2(n98), .B1(B[30]), .B2(n99), .ZN(RES[30]) );
  INV_X1 U82 ( .A(B[30]), .ZN(n98) );
  AOI22_X1 U83 ( .A1(n31), .A2(n100), .B1(A[30]), .B2(n37), .ZN(n97) );
  AOI22_X1 U84 ( .A1(n28), .A2(n100), .B1(A[30]), .B2(n34), .ZN(n99) );
  OAI22_X1 U85 ( .A1(n165), .A2(n166), .B1(B[15]), .B2(n167), .ZN(RES[15]) );
  INV_X1 U86 ( .A(B[15]), .ZN(n166) );
  AOI22_X1 U87 ( .A1(n30), .A2(n1), .B1(A[15]), .B2(n36), .ZN(n165) );
  AOI22_X1 U88 ( .A1(n27), .A2(n1), .B1(A[15]), .B2(n33), .ZN(n167) );
  OAI22_X1 U89 ( .A1(n69), .A2(n70), .B1(B[8]), .B2(n71), .ZN(RES[8]) );
  INV_X1 U90 ( .A(B[8]), .ZN(n70) );
  AOI22_X1 U91 ( .A1(n32), .A2(n20), .B1(A[8]), .B2(n38), .ZN(n69) );
  AOI22_X1 U92 ( .A1(n29), .A2(n20), .B1(A[8]), .B2(n35), .ZN(n71) );
  OAI22_X1 U93 ( .A1(n169), .A2(n170), .B1(B[14]), .B2(n171), .ZN(RES[14]) );
  INV_X1 U94 ( .A(B[14]), .ZN(n170) );
  AOI22_X1 U95 ( .A1(n30), .A2(n26), .B1(A[14]), .B2(n36), .ZN(n169) );
  AOI22_X1 U96 ( .A1(n27), .A2(n26), .B1(A[14]), .B2(n33), .ZN(n171) );
  OAI22_X1 U97 ( .A1(n73), .A2(n8), .B1(B[7]), .B2(n75), .ZN(RES[7]) );
  AOI22_X1 U98 ( .A1(n32), .A2(n19), .B1(A[7]), .B2(n38), .ZN(n73) );
  AOI22_X1 U99 ( .A1(n29), .A2(n19), .B1(A[7]), .B2(n35), .ZN(n75) );
  OAI22_X1 U100 ( .A1(n65), .A2(n9), .B1(B[9]), .B2(n67), .ZN(RES[9]) );
  AOI22_X1 U101 ( .A1(n32), .A2(n21), .B1(n38), .B2(A[9]), .ZN(n65) );
  AOI22_X1 U102 ( .A1(n29), .A2(n21), .B1(n35), .B2(A[9]), .ZN(n67) );
  BUF_X1 U103 ( .A(SEL[0]), .Z(n28) );
  BUF_X1 U104 ( .A(SEL[0]), .Z(n27) );
  BUF_X1 U105 ( .A(SEL[0]), .Z(n29) );
  BUF_X1 U106 ( .A(SEL[1]), .Z(n31) );
  BUF_X1 U107 ( .A(SEL[1]), .Z(n30) );
  BUF_X1 U108 ( .A(SEL[3]), .Z(n37) );
  BUF_X1 U109 ( .A(SEL[2]), .Z(n34) );
  BUF_X1 U110 ( .A(SEL[3]), .Z(n36) );
  BUF_X1 U111 ( .A(SEL[2]), .Z(n33) );
  BUF_X1 U112 ( .A(SEL[1]), .Z(n32) );
  BUF_X1 U113 ( .A(SEL[3]), .Z(n38) );
  BUF_X1 U114 ( .A(SEL[2]), .Z(n35) );
  INV_X1 U115 ( .A(A[15]), .ZN(n1) );
  AOI22_X1 U116 ( .A1(n28), .A2(n136), .B1(A[22]), .B2(n34), .ZN(n135) );
  AOI22_X1 U117 ( .A1(n31), .A2(n136), .B1(A[22]), .B2(n37), .ZN(n133) );
  INV_X1 U118 ( .A(A[22]), .ZN(n136) );
  AOI22_X1 U119 ( .A1(n27), .A2(n160), .B1(A[17]), .B2(n33), .ZN(n159) );
  AOI22_X1 U120 ( .A1(n30), .A2(n160), .B1(A[17]), .B2(n36), .ZN(n157) );
  INV_X1 U121 ( .A(A[17]), .ZN(n160) );
  AOI22_X1 U122 ( .A1(n29), .A2(n16), .B1(A[4]), .B2(n35), .ZN(n87) );
  AOI22_X1 U123 ( .A1(n32), .A2(n16), .B1(A[4]), .B2(n38), .ZN(n85) );
  AOI22_X1 U124 ( .A1(n29), .A2(n18), .B1(A[6]), .B2(n35), .ZN(n79) );
  AOI22_X1 U125 ( .A1(n32), .A2(n18), .B1(A[6]), .B2(n38), .ZN(n77) );
  AOI22_X1 U126 ( .A1(n27), .A2(n13), .B1(A[1]), .B2(n33), .ZN(n147) );
  AOI22_X1 U127 ( .A1(n30), .A2(n13), .B1(A[1]), .B2(n36), .ZN(n145) );
  AOI22_X1 U128 ( .A1(n32), .A2(n17), .B1(A[5]), .B2(n38), .ZN(n81) );
  AOI22_X1 U129 ( .A1(n29), .A2(n17), .B1(A[5]), .B2(n35), .ZN(n83) );
  AOI22_X1 U130 ( .A1(n32), .A2(n15), .B1(A[3]), .B2(n38), .ZN(n89) );
  AOI22_X1 U131 ( .A1(n29), .A2(n15), .B1(A[3]), .B2(n35), .ZN(n91) );
  OAI22_X1 U132 ( .A1(n101), .A2(n4), .B1(B[2]), .B2(n103), .ZN(RES[2]) );
  OAI22_X1 U133 ( .A1(n85), .A2(n6), .B1(B[4]), .B2(n87), .ZN(RES[4]) );
  OAI22_X1 U134 ( .A1(n181), .A2(n10), .B1(B[11]), .B2(n183), .ZN(RES[11]) );
  OAI22_X1 U135 ( .A1(n173), .A2(n11), .B1(B[13]), .B2(n175), .ZN(RES[13]) );
  OAI22_X1 U136 ( .A1(n89), .A2(n5), .B1(B[3]), .B2(n91), .ZN(RES[3]) );
  OAI22_X1 U137 ( .A1(n189), .A2(n2), .B1(B[0]), .B2(n191), .ZN(RES[0]) );
  OAI22_X1 U138 ( .A1(n81), .A2(n7), .B1(B[5]), .B2(n83), .ZN(RES[5]) );
  AOI22_X1 U139 ( .A1(n27), .A2(n12), .B1(A[0]), .B2(n33), .ZN(n191) );
  AOI22_X1 U140 ( .A1(n30), .A2(n12), .B1(A[0]), .B2(n36), .ZN(n189) );
  OAI22_X1 U141 ( .A1(n177), .A2(n178), .B1(B[12]), .B2(n179), .ZN(RES[12]) );
  INV_X1 U142 ( .A(B[12]), .ZN(n178) );
  OAI22_X1 U143 ( .A1(n185), .A2(n186), .B1(B[10]), .B2(n187), .ZN(RES[10]) );
  INV_X1 U144 ( .A(B[10]), .ZN(n186) );
  OAI22_X1 U145 ( .A1(n145), .A2(n3), .B1(B[1]), .B2(n147), .ZN(RES[1]) );
  OAI22_X1 U146 ( .A1(n77), .A2(n78), .B1(B[6]), .B2(n79), .ZN(RES[6]) );
  INV_X1 U147 ( .A(B[6]), .ZN(n78) );
  INV_X1 U148 ( .A(B[0]), .ZN(n2) );
  INV_X1 U149 ( .A(B[1]), .ZN(n3) );
  INV_X1 U150 ( .A(B[2]), .ZN(n4) );
  INV_X1 U151 ( .A(B[3]), .ZN(n5) );
  INV_X1 U152 ( .A(B[4]), .ZN(n6) );
  INV_X1 U153 ( .A(B[5]), .ZN(n7) );
  INV_X1 U154 ( .A(B[7]), .ZN(n8) );
  INV_X1 U155 ( .A(B[9]), .ZN(n9) );
  INV_X1 U156 ( .A(B[11]), .ZN(n10) );
  INV_X1 U157 ( .A(B[13]), .ZN(n11) );
  INV_X1 U158 ( .A(A[0]), .ZN(n12) );
  INV_X1 U159 ( .A(A[1]), .ZN(n13) );
  INV_X1 U160 ( .A(A[2]), .ZN(n14) );
  INV_X1 U161 ( .A(A[3]), .ZN(n15) );
  INV_X1 U162 ( .A(A[4]), .ZN(n16) );
  INV_X1 U163 ( .A(A[5]), .ZN(n17) );
  INV_X1 U164 ( .A(A[6]), .ZN(n18) );
  INV_X1 U165 ( .A(A[7]), .ZN(n19) );
  INV_X1 U166 ( .A(A[8]), .ZN(n20) );
  INV_X1 U167 ( .A(A[9]), .ZN(n21) );
  INV_X1 U168 ( .A(A[10]), .ZN(n22) );
  INV_X1 U169 ( .A(A[11]), .ZN(n23) );
  INV_X1 U170 ( .A(A[12]), .ZN(n24) );
  INV_X1 U171 ( .A(A[13]), .ZN(n25) );
  INV_X1 U172 ( .A(A[14]), .ZN(n26) );
endmodule


module COMPARATOR_NB32_0 ( AdderRes, MSB, CO, OP_CODE, US, SOUT );
  input [31:0] AdderRes;
  input [1:0] MSB;
  input [2:0] OP_CODE;
  output [31:0] SOUT;
  input CO, US;
  wire   n7, n8, n9, n10, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n1, n2;
  assign SOUT[31] = 1'b0;
  assign SOUT[30] = 1'b0;
  assign SOUT[29] = 1'b0;
  assign SOUT[28] = 1'b0;
  assign SOUT[27] = 1'b0;
  assign SOUT[26] = 1'b0;
  assign SOUT[25] = 1'b0;
  assign SOUT[24] = 1'b0;
  assign SOUT[23] = 1'b0;
  assign SOUT[22] = 1'b0;
  assign SOUT[21] = 1'b0;
  assign SOUT[20] = 1'b0;
  assign SOUT[19] = 1'b0;
  assign SOUT[18] = 1'b0;
  assign SOUT[17] = 1'b0;
  assign SOUT[16] = 1'b0;
  assign SOUT[15] = 1'b0;
  assign SOUT[14] = 1'b0;
  assign SOUT[13] = 1'b0;
  assign SOUT[12] = 1'b0;
  assign SOUT[11] = 1'b0;
  assign SOUT[10] = 1'b0;
  assign SOUT[9] = 1'b0;
  assign SOUT[8] = 1'b0;
  assign SOUT[7] = 1'b0;
  assign SOUT[6] = 1'b0;
  assign SOUT[5] = 1'b0;
  assign SOUT[4] = 1'b0;
  assign SOUT[3] = 1'b0;
  assign SOUT[2] = 1'b0;
  assign SOUT[1] = 1'b0;

  NAND3_X1 U28 ( .A1(n1), .A2(n2), .A3(n14), .ZN(n11) );
  NAND3_X1 U29 ( .A1(n15), .A2(n1), .A3(OP_CODE[0]), .ZN(n23) );
  NOR4_X1 U2 ( .A1(AdderRes[9]), .A2(AdderRes[8]), .A3(AdderRes[7]), .A4(
        AdderRes[6]), .ZN(n33) );
  INV_X1 U3 ( .A(n17), .ZN(n15) );
  NOR4_X1 U4 ( .A1(AdderRes[5]), .A2(AdderRes[4]), .A3(AdderRes[3]), .A4(
        AdderRes[31]), .ZN(n32) );
  NOR4_X1 U5 ( .A1(AdderRes[16]), .A2(AdderRes[15]), .A3(AdderRes[14]), .A4(
        AdderRes[13]), .ZN(n27) );
  NOR2_X1 U6 ( .A1(n24), .A2(n25), .ZN(n17) );
  NAND4_X1 U7 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n25) );
  NAND4_X1 U8 ( .A1(n30), .A2(n31), .A3(n32), .A4(n33), .ZN(n24) );
  NOR4_X1 U9 ( .A1(AdderRes[12]), .A2(AdderRes[11]), .A3(AdderRes[10]), .A4(
        AdderRes[0]), .ZN(n26) );
  NOR4_X1 U10 ( .A1(AdderRes[1]), .A2(AdderRes[19]), .A3(AdderRes[18]), .A4(
        AdderRes[17]), .ZN(n28) );
  XNOR2_X1 U11 ( .A(MSB[0]), .B(MSB[1]), .ZN(n20) );
  AOI221_X1 U12 ( .B1(n16), .B2(n17), .C1(CO), .C2(n18), .A(n19), .ZN(n9) );
  NOR3_X1 U13 ( .A1(n2), .A2(OP_CODE[1]), .A3(CO), .ZN(n19) );
  AOI22_X1 U14 ( .A1(MSB[1]), .A2(n21), .B1(MSB[0]), .B2(n18), .ZN(n7) );
  NAND2_X1 U15 ( .A1(n22), .A2(n23), .ZN(n21) );
  INV_X1 U16 ( .A(n16), .ZN(n22) );
  AOI211_X1 U17 ( .C1(OP_CODE[0]), .C2(n17), .A(n2), .B(n1), .ZN(n18) );
  NOR3_X1 U18 ( .A1(OP_CODE[0]), .A2(OP_CODE[1]), .A3(n2), .ZN(n16) );
  OAI221_X1 U19 ( .B1(n7), .B2(n8), .C1(n9), .C2(n10), .A(n11), .ZN(SOUT[0])
         );
  INV_X1 U20 ( .A(n10), .ZN(n8) );
  NOR2_X1 U21 ( .A1(US), .A2(n20), .ZN(n10) );
  XNOR2_X1 U22 ( .A(OP_CODE[0]), .B(n15), .ZN(n14) );
  INV_X1 U23 ( .A(OP_CODE[1]), .ZN(n1) );
  NOR4_X1 U24 ( .A1(AdderRes[30]), .A2(AdderRes[2]), .A3(AdderRes[29]), .A4(
        AdderRes[28]), .ZN(n31) );
  NOR4_X1 U25 ( .A1(AdderRes[23]), .A2(AdderRes[22]), .A3(AdderRes[21]), .A4(
        AdderRes[20]), .ZN(n29) );
  NOR4_X1 U26 ( .A1(AdderRes[27]), .A2(AdderRes[26]), .A3(AdderRes[25]), .A4(
        AdderRes[24]), .ZN(n30) );
  INV_X1 U27 ( .A(OP_CODE[2]), .ZN(n2) );
endmodule


module SHIFTER_NB32_LS5_0 ( FUNC, US, DATA1, DATA2, OUTSHFT );
  input [1:0] FUNC;
  input [31:0] DATA1;
  input [4:0] DATA2;
  output [31:0] OUTSHFT;
  input US;
  wire   n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n344, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n609, n612, n615, n617, n620,
         n622, n624, n626, n627, n628, n629, n630, n631, n632, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n668, n669, n671,
         n672, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39;

  NOR2_X2 U548 ( .A1(n242), .A2(n21), .ZN(n154) );
  NOR2_X2 U551 ( .A1(n241), .A2(n21), .ZN(n152) );
  NAND3_X1 U619 ( .A1(n140), .A2(n141), .A3(n142), .ZN(OUTSHFT[9]) );
  NAND3_X1 U620 ( .A1(n158), .A2(n159), .A3(n160), .ZN(OUTSHFT[8]) );
  NAND3_X1 U621 ( .A1(n168), .A2(n169), .A3(n170), .ZN(OUTSHFT[7]) );
  NAND3_X1 U622 ( .A1(n179), .A2(n180), .A3(n181), .ZN(OUTSHFT[6]) );
  NAND3_X1 U623 ( .A1(n190), .A2(n191), .A3(n192), .ZN(OUTSHFT[5]) );
  NAND3_X1 U624 ( .A1(n201), .A2(n202), .A3(n203), .ZN(OUTSHFT[4]) );
  NAND3_X1 U625 ( .A1(n303), .A2(n304), .A3(n305), .ZN(OUTSHFT[27]) );
  NAND3_X1 U626 ( .A1(n468), .A2(n20), .A3(n312), .ZN(n467) );
  NAND3_X1 U627 ( .A1(n559), .A2(n560), .A3(n561), .ZN(OUTSHFT[14]) );
  NAND3_X1 U628 ( .A1(n571), .A2(n572), .A3(n573), .ZN(OUTSHFT[13]) );
  NAND3_X1 U629 ( .A1(n643), .A2(n644), .A3(n645), .ZN(OUTSHFT[11]) );
  NAND3_X1 U630 ( .A1(n678), .A2(n679), .A3(n680), .ZN(OUTSHFT[10]) );
  NAND2_X2 U2 ( .A1(DATA2[2]), .A2(n20), .ZN(n339) );
  NAND2_X2 U3 ( .A1(n19), .A2(n20), .ZN(n341) );
  INV_X2 U4 ( .A(n13), .ZN(n14) );
  INV_X2 U5 ( .A(n353), .ZN(n12) );
  NAND2_X2 U6 ( .A1(DATA2[2]), .A2(DATA2[3]), .ZN(n353) );
  INV_X2 U7 ( .A(n336), .ZN(n16) );
  INV_X2 U8 ( .A(n546), .ZN(n156) );
  BUF_X2 U9 ( .A(n143), .Z(n17) );
  INV_X2 U10 ( .A(n11), .ZN(n10) );
  INV_X2 U11 ( .A(n6), .ZN(n5) );
  INV_X4 U12 ( .A(n1), .ZN(n4) );
  AOI222_X1 U13 ( .A1(n5), .A2(DATA1[1]), .B1(n11), .B2(DATA1[0]), .C1(n4), 
        .C2(n25), .ZN(n268) );
  NOR2_X1 U14 ( .A1(n241), .A2(n22), .ZN(n312) );
  OR2_X1 U15 ( .A1(DATA2[0]), .A2(DATA2[1]), .ZN(n1) );
  OAI21_X1 U16 ( .B1(n437), .B2(n353), .A(n566), .ZN(n252) );
  INV_X1 U17 ( .A(n640), .ZN(n383) );
  INV_X1 U18 ( .A(n658), .ZN(n313) );
  INV_X1 U19 ( .A(n358), .ZN(n456) );
  INV_X1 U20 ( .A(n490), .ZN(n487) );
  INV_X1 U21 ( .A(n271), .ZN(n267) );
  INV_X1 U22 ( .A(n395), .ZN(n176) );
  AOI222_X1 U23 ( .A1(n413), .A2(n15), .B1(n414), .B2(n16), .C1(n399), .C2(n14), .ZN(n658) );
  AOI222_X1 U24 ( .A1(n362), .A2(n15), .B1(n363), .B2(n16), .C1(n344), .C2(n14), .ZN(n595) );
  AOI222_X1 U25 ( .A1(n425), .A2(n15), .B1(n441), .B2(n16), .C1(n426), .C2(n14), .ZN(n566) );
  AOI211_X1 U26 ( .C1(n637), .C2(n12), .A(n638), .B(n639), .ZN(n291) );
  OAI22_X1 U27 ( .A1(n336), .A2(n382), .B1(n339), .B2(n383), .ZN(n639) );
  INV_X1 U28 ( .A(n311), .ZN(n292) );
  OAI221_X1 U29 ( .B1(n552), .B2(n339), .C1(n500), .C2(n341), .A(n553), .ZN(
        n244) );
  INV_X1 U30 ( .A(n399), .ZN(n552) );
  AOI22_X1 U31 ( .A1(n12), .A2(n414), .B1(n16), .B2(n413), .ZN(n553) );
  OAI221_X1 U32 ( .B1(n432), .B2(n339), .C1(n433), .C2(n341), .A(n570), .ZN(
        n257) );
  AOI22_X1 U33 ( .A1(n12), .A2(n520), .B1(n16), .B2(n521), .ZN(n570) );
  OAI221_X1 U34 ( .B1(n500), .B2(n339), .C1(n396), .C2(n341), .A(n501), .ZN(
        n223) );
  AOI22_X1 U35 ( .A1(n12), .A2(n413), .B1(n16), .B2(n399), .ZN(n501) );
  OAI221_X1 U36 ( .B1(n352), .B2(n339), .C1(n455), .C2(n341), .A(n533), .ZN(
        n490) );
  AOI22_X1 U37 ( .A1(n12), .A2(n453), .B1(n16), .B2(n454), .ZN(n533) );
  OAI221_X1 U38 ( .B1(n428), .B2(n339), .C1(n432), .C2(n341), .A(n519), .ZN(
        n271) );
  AOI22_X1 U39 ( .A1(n12), .A2(n431), .B1(n16), .B2(n520), .ZN(n519) );
  OAI221_X1 U40 ( .B1(n531), .B2(n339), .C1(n449), .C2(n341), .A(n532), .ZN(
        n488) );
  INV_X1 U41 ( .A(n344), .ZN(n531) );
  AOI22_X1 U42 ( .A1(n12), .A2(n363), .B1(n16), .B2(n362), .ZN(n532) );
  OAI221_X1 U43 ( .B1(n360), .B2(n353), .C1(n361), .C2(n336), .A(n337), .ZN(
        n155) );
  OAI221_X1 U44 ( .B1(n523), .B2(n353), .C1(n437), .C2(n336), .A(n691), .ZN(
        n327) );
  OAI221_X1 U45 ( .B1(n455), .B2(n339), .C1(n456), .C2(n341), .A(n606), .ZN(
        n282) );
  AOI22_X1 U46 ( .A1(n12), .A2(n454), .B1(n16), .B2(n534), .ZN(n606) );
  OAI221_X1 U47 ( .B1(n470), .B2(n339), .C1(n372), .C2(n341), .A(n471), .ZN(
        n204) );
  AOI22_X1 U48 ( .A1(n12), .A2(n389), .B1(n16), .B2(n375), .ZN(n471) );
  OAI221_X1 U49 ( .B1(n401), .B2(n353), .C1(n402), .C2(n336), .A(n557), .ZN(
        n239) );
  AOI22_X1 U50 ( .A1(n15), .A2(n558), .B1(n14), .B2(n506), .ZN(n557) );
  OAI221_X1 U51 ( .B1(n449), .B2(n339), .C1(n338), .C2(n341), .A(n450), .ZN(
        n193) );
  AOI22_X1 U52 ( .A1(n12), .A2(n362), .B1(n16), .B2(n344), .ZN(n450) );
  OAI221_X1 U53 ( .B1(n8), .B2(n27), .C1(n6), .C2(n24), .A(n726), .ZN(n640) );
  AOI21_X1 U54 ( .B1(n25), .B2(n11), .A(n541), .ZN(n726) );
  OAI221_X1 U55 ( .B1(n712), .B2(n339), .C1(n470), .C2(n341), .A(n713), .ZN(
        n539) );
  INV_X1 U56 ( .A(n375), .ZN(n712) );
  AOI22_X1 U57 ( .A1(n12), .A2(n390), .B1(n16), .B2(n389), .ZN(n713) );
  OAI221_X1 U58 ( .B1(n396), .B2(n339), .C1(n397), .C2(n341), .A(n398), .ZN(
        n171) );
  AOI22_X1 U59 ( .A1(n12), .A2(n399), .B1(n16), .B2(n400), .ZN(n398) );
  OAI221_X1 U60 ( .B1(n455), .B2(n353), .C1(n456), .C2(n336), .A(n457), .ZN(
        n200) );
  OAI221_X1 U61 ( .B1(n432), .B2(n353), .C1(n433), .C2(n336), .A(n434), .ZN(
        n189) );
  OAI221_X1 U62 ( .B1(n406), .B2(n353), .C1(n407), .C2(n336), .A(n408), .ZN(
        n178) );
  OAI221_X1 U63 ( .B1(n382), .B2(n353), .C1(n383), .C2(n336), .A(n384), .ZN(
        n167) );
  OAI221_X1 U64 ( .B1(n432), .B2(n336), .C1(n433), .C2(n339), .A(n698), .ZN(
        n321) );
  AOI21_X1 U65 ( .B1(n12), .B2(n521), .A(n699), .ZN(n698) );
  INV_X1 U66 ( .A(n683), .ZN(n699) );
  OAI221_X1 U67 ( .B1(n377), .B2(n353), .C1(n378), .C2(n336), .A(n725), .ZN(
        n543) );
  AOI22_X1 U68 ( .A1(n15), .A2(n641), .B1(n14), .B2(n640), .ZN(n725) );
  INV_X1 U69 ( .A(n466), .ZN(n314) );
  OAI22_X1 U70 ( .A1(n448), .A2(n341), .B1(n335), .B2(n339), .ZN(n198) );
  OAI22_X1 U71 ( .A1(n421), .A2(n341), .B1(n268), .B2(n339), .ZN(n187) );
  NAND2_X1 U72 ( .A1(n152), .A2(n14), .ZN(n221) );
  AOI22_X1 U73 ( .A1(n413), .A2(n14), .B1(n414), .B2(n15), .ZN(n395) );
  OAI22_X1 U74 ( .A1(n466), .A2(n530), .B1(n335), .B2(n499), .ZN(n529) );
  INV_X1 U75 ( .A(n488), .ZN(n530) );
  AOI22_X1 U76 ( .A1(n389), .A2(n14), .B1(n390), .B2(n15), .ZN(n371) );
  AOI22_X1 U77 ( .A1(n362), .A2(n14), .B1(n363), .B2(n15), .ZN(n337) );
  AOI22_X1 U78 ( .A1(n425), .A2(n14), .B1(n441), .B2(n15), .ZN(n691) );
  AOI22_X1 U79 ( .A1(n375), .A2(n14), .B1(n389), .B2(n15), .ZN(n632) );
  OAI21_X1 U80 ( .B1(n335), .B2(n353), .A(n595), .ZN(n285) );
  OAI21_X1 U81 ( .B1(n335), .B2(n336), .A(n337), .ZN(n153) );
  OAI22_X1 U82 ( .A1(n516), .A2(n466), .B1(n268), .B2(n499), .ZN(n515) );
  INV_X1 U83 ( .A(n269), .ZN(n516) );
  OAI22_X1 U84 ( .A1(n498), .A2(n466), .B1(n220), .B2(n499), .ZN(n497) );
  INV_X1 U85 ( .A(n223), .ZN(n498) );
  NAND2_X1 U86 ( .A1(n312), .A2(n14), .ZN(n499) );
  OAI21_X1 U87 ( .B1(n280), .B2(n339), .A(n354), .ZN(n146) );
  OAI21_X1 U88 ( .B1(n254), .B2(n339), .A(n683), .ZN(n328) );
  AOI21_X1 U89 ( .B1(n299), .B2(n415), .A(n292), .ZN(n365) );
  INV_X1 U90 ( .A(n174), .ZN(n415) );
  OAI211_X1 U91 ( .C1(n352), .C2(n353), .A(n354), .B(n355), .ZN(n157) );
  AOI22_X1 U92 ( .A1(n16), .A2(n356), .B1(n15), .B2(n358), .ZN(n355) );
  NOR3_X1 U93 ( .A1(n341), .A2(n311), .A3(n1), .ZN(n549) );
  OAI21_X1 U94 ( .B1(n254), .B2(n336), .A(n434), .ZN(n183) );
  BUF_X1 U95 ( .A(n581), .Z(n7) );
  OAI21_X1 U96 ( .B1(n254), .B2(n353), .A(n522), .ZN(n272) );
  BUF_X1 U97 ( .A(n581), .Z(n8) );
  BUF_X1 U98 ( .A(n581), .Z(n9) );
  OAI21_X1 U99 ( .B1(n442), .B2(n339), .A(n174), .ZN(n329) );
  OAI21_X1 U100 ( .B1(n280), .B2(n336), .A(n457), .ZN(n194) );
  AOI22_X1 U101 ( .A1(n302), .A2(n21), .B1(n22), .B2(n288), .ZN(n301) );
  OAI21_X1 U102 ( .B1(n280), .B2(n353), .A(n535), .ZN(n491) );
  OAI21_X1 U103 ( .B1(n336), .B2(n234), .A(n408), .ZN(n172) );
  OAI21_X1 U104 ( .B1(n361), .B2(n353), .A(n595), .ZN(n278) );
  OAI21_X1 U105 ( .B1(n442), .B2(n353), .A(n522), .ZN(n273) );
  OAI21_X1 U106 ( .B1(n7), .B2(n23), .A(n280), .ZN(n358) );
  OAI21_X1 U107 ( .B1(n336), .B2(n370), .A(n371), .ZN(n165) );
  OAI21_X1 U108 ( .B1(n456), .B2(n353), .A(n535), .ZN(n485) );
  OAI21_X1 U109 ( .B1(n433), .B2(n353), .A(n522), .ZN(n265) );
  OAI21_X1 U110 ( .B1(n407), .B2(n353), .A(n505), .ZN(n216) );
  OAI21_X1 U111 ( .B1(n268), .B2(n353), .A(n566), .ZN(n260) );
  OAI21_X1 U112 ( .B1(n383), .B2(n353), .A(n475), .ZN(n212) );
  OAI21_X1 U113 ( .B1(n268), .B2(n336), .A(n691), .ZN(n326) );
  AOI22_X1 U114 ( .A1(n171), .A2(n314), .B1(n176), .B2(n312), .ZN(n394) );
  AOI22_X1 U115 ( .A1(n161), .A2(n314), .B1(n165), .B2(n312), .ZN(n369) );
  AOI22_X1 U116 ( .A1(n285), .A2(n21), .B1(n22), .B2(n283), .ZN(n284) );
  NOR2_X1 U117 ( .A1(n341), .A2(n297), .ZN(n638) );
  OAI21_X1 U118 ( .B1(n442), .B2(n336), .A(n207), .ZN(n185) );
  NAND2_X1 U119 ( .A1(n299), .A2(n14), .ZN(n235) );
  NAND2_X1 U120 ( .A1(DATA2[3]), .A2(n19), .ZN(n336) );
  INV_X1 U121 ( .A(n339), .ZN(n15) );
  INV_X1 U122 ( .A(n702), .ZN(n433) );
  OAI221_X1 U123 ( .B1(n10), .B2(n23), .C1(n7), .C2(n24), .A(n254), .ZN(n702)
         );
  INV_X1 U124 ( .A(n707), .ZN(n437) );
  OAI21_X1 U125 ( .B1(n233), .B2(n8), .A(n268), .ZN(n707) );
  INV_X1 U126 ( .A(n414), .ZN(n220) );
  INV_X1 U127 ( .A(n370), .ZN(n541) );
  NOR2_X1 U128 ( .A1(DATA2[3]), .A2(n310), .ZN(n646) );
  INV_X1 U129 ( .A(n356), .ZN(n455) );
  INV_X1 U130 ( .A(n504), .ZN(n401) );
  INV_X1 U131 ( .A(n474), .ZN(n377) );
  NOR2_X1 U132 ( .A1(DATA2[3]), .A2(n210), .ZN(n208) );
  INV_X1 U133 ( .A(n641), .ZN(n382) );
  INV_X1 U134 ( .A(n558), .ZN(n406) );
  INV_X1 U135 ( .A(n534), .ZN(n352) );
  INV_X1 U136 ( .A(n637), .ZN(n378) );
  INV_X1 U137 ( .A(n475), .ZN(n205) );
  INV_X1 U138 ( .A(n363), .ZN(n448) );
  INV_X1 U139 ( .A(n441), .ZN(n421) );
  INV_X1 U140 ( .A(n390), .ZN(n476) );
  NAND2_X1 U141 ( .A1(n505), .A2(n207), .ZN(n229) );
  BUF_X1 U142 ( .A(n341), .Z(n13) );
  INV_X1 U143 ( .A(n426), .ZN(n517) );
  INV_X1 U144 ( .A(n431), .ZN(n568) );
  INV_X1 U145 ( .A(n521), .ZN(n428) );
  INV_X1 U146 ( .A(n400), .ZN(n500) );
  INV_X1 U147 ( .A(n454), .ZN(n348) );
  INV_X1 U148 ( .A(n520), .ZN(n427) );
  INV_X1 U149 ( .A(n453), .ZN(n347) );
  INV_X1 U150 ( .A(n506), .ZN(n407) );
  INV_X1 U151 ( .A(n227), .ZN(n218) );
  INV_X1 U152 ( .A(n384), .ZN(n162) );
  INV_X1 U153 ( .A(n468), .ZN(n210) );
  INV_X1 U154 ( .A(n234), .ZN(n648) );
  INV_X1 U155 ( .A(n564), .ZN(n255) );
  OAI21_X1 U156 ( .B1(n442), .B2(n341), .A(n298), .ZN(n564) );
  INV_X1 U157 ( .A(n207), .ZN(n480) );
  INV_X1 U158 ( .A(n447), .ZN(n446) );
  AOI22_X1 U159 ( .A1(n193), .A2(n314), .B1(n198), .B2(n312), .ZN(n447) );
  INV_X1 U160 ( .A(n420), .ZN(n419) );
  AOI22_X1 U161 ( .A1(n182), .A2(n314), .B1(n187), .B2(n312), .ZN(n420) );
  INV_X1 U162 ( .A(n334), .ZN(n333) );
  AOI22_X1 U163 ( .A1(n144), .A2(n314), .B1(n153), .B2(n312), .ZN(n334) );
  INV_X1 U164 ( .A(n324), .ZN(n323) );
  AOI22_X1 U165 ( .A1(n314), .A2(n325), .B1(n326), .B2(n312), .ZN(n324) );
  AOI222_X1 U166 ( .A1(n350), .A2(n15), .B1(n359), .B2(n16), .C1(n351), .C2(
        n14), .ZN(n535) );
  AOI222_X1 U167 ( .A1(n435), .A2(n15), .B1(n436), .B2(n16), .C1(n430), .C2(
        n14), .ZN(n522) );
  AOI21_X1 U168 ( .B1(n3), .B2(n5), .A(n682), .ZN(n254) );
  OAI221_X1 U169 ( .B1(n10), .B2(n34), .C1(n7), .C2(n33), .A(n717), .ZN(n375)
         );
  AOI22_X1 U170 ( .A1(DATA1[11]), .A2(n5), .B1(DATA1[12]), .B2(n4), .ZN(n717)
         );
  AOI21_X1 U171 ( .B1(n3), .B2(n11), .A(n577), .ZN(n280) );
  NAND2_X1 U172 ( .A1(n219), .A2(n309), .ZN(n150) );
  OAI221_X1 U173 ( .B1(n579), .B2(n29), .C1(n8), .C2(n28), .A(n675), .ZN(n413)
         );
  OAI221_X1 U174 ( .B1(n10), .B2(n31), .C1(n8), .C2(n30), .A(n626), .ZN(n362)
         );
  AOI22_X1 U175 ( .A1(DATA1[8]), .A2(n5), .B1(DATA1[9]), .B2(n4), .ZN(n626) );
  OAI221_X1 U176 ( .B1(n10), .B2(n32), .C1(n7), .C2(n31), .A(n706), .ZN(n425)
         );
  AOI22_X1 U177 ( .A1(DATA1[9]), .A2(n5), .B1(DATA1[10]), .B2(n4), .ZN(n706)
         );
  OAI221_X1 U178 ( .B1(n10), .B2(n33), .C1(n581), .C2(n32), .A(n672), .ZN(n399) );
  AOI22_X1 U179 ( .A1(DATA1[10]), .A2(n5), .B1(DATA1[11]), .B2(n4), .ZN(n672)
         );
  OAI221_X1 U180 ( .B1(n579), .B2(n35), .C1(n9), .C2(n34), .A(n622), .ZN(n344)
         );
  AOI22_X1 U181 ( .A1(DATA1[12]), .A2(n5), .B1(DATA1[13]), .B2(n4), .ZN(n622)
         );
  OAI221_X1 U182 ( .B1(n10), .B2(n30), .C1(n8), .C2(n29), .A(n714), .ZN(n389)
         );
  AOI22_X1 U183 ( .A1(DATA1[7]), .A2(n5), .B1(DATA1[8]), .B2(n4), .ZN(n714) );
  OAI221_X1 U184 ( .B1(n10), .B2(n24), .C1(n581), .C2(n23), .A(n674), .ZN(n414) );
  OAI221_X1 U185 ( .B1(n10), .B2(n27), .C1(n8), .C2(n26), .A(n624), .ZN(n363)
         );
  OAI221_X1 U186 ( .B1(n10), .B2(n28), .C1(n7), .C2(n27), .A(n705), .ZN(n441)
         );
  INV_X1 U187 ( .A(n219), .ZN(n238) );
  AOI222_X1 U188 ( .A1(n385), .A2(n15), .B1(n386), .B2(n16), .C1(n380), .C2(
        n14), .ZN(n475) );
  INV_X1 U189 ( .A(n173), .ZN(n145) );
  OAI221_X1 U190 ( .B1(n340), .B2(n339), .C1(n360), .C2(n341), .A(n578), .ZN(
        n283) );
  AOI22_X1 U191 ( .A1(n12), .A2(n346), .B1(n16), .B2(n451), .ZN(n578) );
  OAI221_X1 U192 ( .B1(n422), .B2(n353), .C1(n423), .C2(n336), .A(n565), .ZN(
        n258) );
  AOI22_X1 U193 ( .A1(n15), .A2(n439), .B1(n14), .B2(n440), .ZN(n565) );
  OAI221_X1 U194 ( .B1(n10), .B2(n602), .C1(n7), .C2(n650), .A(n697), .ZN(n431) );
  AOI22_X1 U195 ( .A1(DATA1[15]), .A2(n5), .B1(DATA1[14]), .B2(n4), .ZN(n697)
         );
  OAI221_X1 U196 ( .B1(n10), .B2(n32), .C1(n7), .C2(n33), .A(n701), .ZN(n521)
         );
  OAI221_X1 U197 ( .B1(n10), .B2(n37), .C1(n8), .C2(n36), .A(n653), .ZN(n400)
         );
  AOI22_X1 U198 ( .A1(DATA1[14]), .A2(n5), .B1(DATA1[15]), .B2(n4), .ZN(n653)
         );
  OAI221_X1 U199 ( .B1(n10), .B2(n2), .C1(n9), .C2(n602), .A(n603), .ZN(n453)
         );
  AOI22_X1 U200 ( .A1(DATA1[14]), .A2(n584), .B1(DATA1[13]), .B2(n4), .ZN(n603) );
  OAI221_X1 U201 ( .B1(n10), .B2(n35), .C1(n9), .C2(n36), .A(n612), .ZN(n454)
         );
  AOI22_X1 U202 ( .A1(DATA1[10]), .A2(n584), .B1(DATA1[9]), .B2(n4), .ZN(n612)
         );
  OAI221_X1 U203 ( .B1(n579), .B2(n36), .C1(n581), .C2(n37), .A(n696), .ZN(
        n520) );
  AOI22_X1 U204 ( .A1(DATA1[11]), .A2(n5), .B1(DATA1[10]), .B2(n4), .ZN(n696)
         );
  OAI221_X1 U205 ( .B1(n8), .B2(n26), .C1(n6), .C2(n23), .A(n666), .ZN(n506)
         );
  OAI221_X1 U206 ( .B1(n373), .B2(n339), .C1(n387), .C2(n341), .A(n642), .ZN(
        n288) );
  AOI22_X1 U207 ( .A1(n12), .A2(n376), .B1(n16), .B2(n472), .ZN(n642) );
  OAI221_X1 U208 ( .B1(n10), .B2(n26), .C1(n7), .C2(n24), .A(n715), .ZN(n390)
         );
  OAI221_X1 U209 ( .B1(n10), .B2(n36), .C1(n581), .C2(n35), .A(n688), .ZN(n426) );
  AOI22_X1 U210 ( .A1(DATA1[13]), .A2(n5), .B1(DATA1[14]), .B2(n4), .ZN(n688)
         );
  NOR2_X1 U211 ( .A1(n154), .A2(n152), .ZN(n466) );
  OAI221_X1 U212 ( .B1(n388), .B2(n339), .C1(n476), .C2(n341), .A(n477), .ZN(
        n211) );
  AOI22_X1 U213 ( .A1(n12), .A2(n478), .B1(n16), .B2(n479), .ZN(n477) );
  OAI221_X1 U214 ( .B1(n361), .B2(n339), .C1(n448), .C2(n341), .A(n458), .ZN(
        n199) );
  AOI22_X1 U215 ( .A1(n12), .A2(n459), .B1(n16), .B2(n460), .ZN(n458) );
  OAI221_X1 U216 ( .B1(n437), .B2(n339), .C1(n421), .C2(n341), .A(n438), .ZN(
        n188) );
  AOI22_X1 U217 ( .A1(n12), .A2(n439), .B1(n16), .B2(n440), .ZN(n438) );
  OAI221_X1 U218 ( .B1(n347), .B2(n339), .C1(n348), .C2(n341), .A(n349), .ZN(
        n151) );
  AOI22_X1 U219 ( .A1(n12), .A2(n350), .B1(n16), .B2(n351), .ZN(n349) );
  OAI221_X1 U220 ( .B1(n402), .B2(n339), .C1(n406), .C2(n341), .A(n503), .ZN(
        n227) );
  AOI22_X1 U221 ( .A1(n12), .A2(n405), .B1(n16), .B2(n504), .ZN(n503) );
  INV_X1 U222 ( .A(n309), .ZN(n299) );
  OAI221_X1 U223 ( .B1(n517), .B2(n339), .C1(n422), .C2(n341), .A(n518), .ZN(
        n269) );
  AOI22_X1 U224 ( .A1(n12), .A2(n441), .B1(n16), .B2(n425), .ZN(n518) );
  OAI221_X1 U225 ( .B1(n348), .B2(n339), .C1(n352), .C2(n341), .A(n452), .ZN(
        n197) );
  AOI22_X1 U226 ( .A1(n12), .A2(n351), .B1(n16), .B2(n453), .ZN(n452) );
  OAI221_X1 U227 ( .B1(n427), .B2(n339), .C1(n428), .C2(n341), .A(n429), .ZN(
        n186) );
  AOI22_X1 U228 ( .A1(n12), .A2(n430), .B1(n16), .B2(n431), .ZN(n429) );
  OAI221_X1 U229 ( .B1(n401), .B2(n339), .C1(n402), .C2(n341), .A(n403), .ZN(
        n175) );
  AOI22_X1 U230 ( .A1(n12), .A2(n404), .B1(n16), .B2(n405), .ZN(n403) );
  OAI221_X1 U231 ( .B1(n360), .B2(n339), .C1(n361), .C2(n341), .A(n536), .ZN(
        n484) );
  AOI22_X1 U232 ( .A1(n12), .A2(n451), .B1(n16), .B2(n459), .ZN(n536) );
  OAI221_X1 U233 ( .B1(n523), .B2(n339), .C1(n437), .C2(n341), .A(n524), .ZN(
        n264) );
  AOI22_X1 U234 ( .A1(n12), .A2(n525), .B1(n16), .B2(n439), .ZN(n524) );
  OAI221_X1 U235 ( .B1(n412), .B2(n339), .C1(n220), .C2(n341), .A(n508), .ZN(
        n215) );
  AOI22_X1 U236 ( .A1(n12), .A2(n509), .B1(n16), .B2(n510), .ZN(n508) );
  OAI221_X1 U237 ( .B1(n411), .B2(n353), .C1(n412), .C2(n336), .A(n395), .ZN(
        n177) );
  OAI221_X1 U238 ( .B1(n387), .B2(n353), .C1(n388), .C2(n336), .A(n371), .ZN(
        n166) );
  OAI221_X1 U239 ( .B1(n377), .B2(n339), .C1(n378), .C2(n341), .A(n379), .ZN(
        n164) );
  AOI22_X1 U240 ( .A1(n12), .A2(n380), .B1(n16), .B2(n381), .ZN(n379) );
  OAI221_X1 U241 ( .B1(n387), .B2(n339), .C1(n388), .C2(n341), .A(n718), .ZN(
        n544) );
  AOI22_X1 U242 ( .A1(n12), .A2(n472), .B1(n16), .B2(n478), .ZN(n718) );
  OAI221_X1 U243 ( .B1(n402), .B2(n353), .C1(n406), .C2(n336), .A(n664), .ZN(
        n316) );
  AOI22_X1 U244 ( .A1(n15), .A2(n506), .B1(n14), .B2(n410), .ZN(n664) );
  OAI221_X1 U245 ( .B1(n411), .B2(n339), .C1(n412), .C2(n341), .A(n551), .ZN(
        n245) );
  AOI22_X1 U246 ( .A1(n12), .A2(n502), .B1(n16), .B2(n509), .ZN(n551) );
  OAI221_X1 U247 ( .B1(n378), .B2(n339), .C1(n382), .C2(n341), .A(n473), .ZN(
        n209) );
  AOI22_X1 U248 ( .A1(n12), .A2(n381), .B1(n16), .B2(n474), .ZN(n473) );
  OAI221_X1 U249 ( .B1(n730), .B2(n339), .C1(n634), .C2(n341), .A(n731), .ZN(
        n542) );
  INV_X1 U250 ( .A(n380), .ZN(n730) );
  AOI22_X1 U251 ( .A1(n12), .A2(n386), .B1(n16), .B2(n385), .ZN(n731) );
  AOI21_X1 U252 ( .B1(n1), .B2(n3), .A(n682), .ZN(n442) );
  OAI221_X1 U253 ( .B1(n579), .B2(n27), .C1(n9), .C2(n28), .A(n620), .ZN(n356)
         );
  OAI221_X1 U254 ( .B1(n10), .B2(n29), .C1(n581), .C2(n30), .A(n668), .ZN(n558) );
  OAI221_X1 U255 ( .B1(n579), .B2(n30), .C1(n581), .C2(n31), .A(n727), .ZN(
        n641) );
  OAI221_X1 U256 ( .B1(n10), .B2(n31), .C1(n9), .C2(n32), .A(n609), .ZN(n534)
         );
  OAI221_X1 U257 ( .B1(n10), .B2(n37), .C1(n8), .C2(n38), .A(n662), .ZN(n504)
         );
  AOI22_X1 U258 ( .A1(DATA1[12]), .A2(n5), .B1(DATA1[11]), .B2(n4), .ZN(n662)
         );
  OAI221_X1 U259 ( .B1(n579), .B2(n38), .C1(n581), .C2(n2), .A(n729), .ZN(n474) );
  AOI22_X1 U260 ( .A1(DATA1[13]), .A2(n5), .B1(DATA1[12]), .B2(n4), .ZN(n729)
         );
  OAI221_X1 U261 ( .B1(n422), .B2(n339), .C1(n423), .C2(n341), .A(n424), .ZN(
        n182) );
  AOI22_X1 U262 ( .A1(n12), .A2(n425), .B1(n16), .B2(n426), .ZN(n424) );
  OAI221_X1 U263 ( .B1(n338), .B2(n339), .C1(n340), .C2(n341), .A(n342), .ZN(
        n144) );
  AOI22_X1 U264 ( .A1(n12), .A2(n344), .B1(n16), .B2(n346), .ZN(n342) );
  OAI221_X1 U265 ( .B1(n567), .B2(n339), .C1(n568), .C2(n341), .A(n569), .ZN(
        n251) );
  INV_X1 U266 ( .A(n430), .ZN(n567) );
  AOI22_X1 U267 ( .A1(n12), .A2(n436), .B1(n16), .B2(n435), .ZN(n569) );
  OAI221_X1 U268 ( .B1(n554), .B2(n339), .C1(n555), .C2(n341), .A(n556), .ZN(
        n237) );
  INV_X1 U269 ( .A(n404), .ZN(n554) );
  AOI22_X1 U270 ( .A1(n12), .A2(n410), .B1(n16), .B2(n409), .ZN(n556) );
  OAI221_X1 U271 ( .B1(n568), .B2(n339), .C1(n427), .C2(n341), .A(n693), .ZN(
        n322) );
  AOI22_X1 U272 ( .A1(n12), .A2(n435), .B1(n16), .B2(n430), .ZN(n693) );
  OAI221_X1 U273 ( .B1(n634), .B2(n339), .C1(n377), .C2(n341), .A(n635), .ZN(
        n289) );
  AOI22_X1 U274 ( .A1(n12), .A2(n385), .B1(n16), .B2(n380), .ZN(n635) );
  OAI221_X1 U275 ( .B1(n388), .B2(n353), .C1(n476), .C2(n336), .A(n632), .ZN(
        n293) );
  OAI221_X1 U276 ( .B1(n555), .B2(n339), .C1(n401), .C2(n341), .A(n659), .ZN(
        n317) );
  AOI22_X1 U277 ( .A1(n12), .A2(n409), .B1(n16), .B2(n404), .ZN(n659) );
  OAI221_X1 U278 ( .B1(n397), .B2(n339), .C1(n411), .C2(n341), .A(n649), .ZN(
        n315) );
  AOI22_X1 U279 ( .A1(n12), .A2(n400), .B1(n16), .B2(n502), .ZN(n649) );
  OAI221_X1 U280 ( .B1(n372), .B2(n339), .C1(n373), .C2(n341), .A(n374), .ZN(
        n161) );
  AOI22_X1 U281 ( .A1(n12), .A2(n375), .B1(n16), .B2(n376), .ZN(n374) );
  OAI221_X1 U282 ( .B1(n579), .B2(n34), .C1(n581), .C2(n35), .A(n728), .ZN(
        n637) );
  AOI22_X1 U283 ( .A1(DATA1[9]), .A2(n5), .B1(DATA1[8]), .B2(n4), .ZN(n728) );
  OAI221_X1 U284 ( .B1(n596), .B2(n339), .C1(n347), .C2(n341), .A(n597), .ZN(
        n277) );
  INV_X1 U285 ( .A(n351), .ZN(n596) );
  AOI22_X1 U286 ( .A1(n12), .A2(n359), .B1(n16), .B2(n350), .ZN(n597) );
  AOI221_X1 U287 ( .B1(n156), .B2(n251), .C1(n17), .C2(n252), .A(n253), .ZN(
        n250) );
  OAI22_X1 U288 ( .A1(n254), .A2(n235), .B1(n255), .B2(n256), .ZN(n253) );
  AOI22_X1 U289 ( .A1(n238), .A2(n257), .B1(n154), .B2(n258), .ZN(n249) );
  AOI22_X1 U290 ( .A1(n154), .A2(n293), .B1(n156), .B2(n636), .ZN(n630) );
  INV_X1 U291 ( .A(n291), .ZN(n636) );
  OAI22_X1 U292 ( .A1(n1), .A2(n615), .B1(n6), .B2(n617), .ZN(n577) );
  AOI22_X1 U293 ( .A1(n385), .A2(n14), .B1(n386), .B2(n15), .ZN(n384) );
  OAI22_X1 U294 ( .A1(n487), .A2(n219), .B1(n335), .B2(n221), .ZN(n486) );
  AOI22_X1 U295 ( .A1(n350), .A2(n14), .B1(n359), .B2(n15), .ZN(n457) );
  AOI22_X1 U296 ( .A1(n435), .A2(n14), .B1(n436), .B2(n15), .ZN(n434) );
  AOI22_X1 U297 ( .A1(n409), .A2(n14), .B1(n410), .B2(n15), .ZN(n408) );
  NOR2_X1 U298 ( .A1(n1), .A2(n617), .ZN(n682) );
  AOI22_X1 U299 ( .A1(n404), .A2(n14), .B1(n409), .B2(n15), .ZN(n507) );
  OAI22_X1 U300 ( .A1(n267), .A2(n219), .B1(n268), .B2(n221), .ZN(n266) );
  OAI22_X1 U301 ( .A1(n218), .A2(n219), .B1(n220), .B2(n221), .ZN(n217) );
  OAI22_X1 U302 ( .A1(n297), .A2(n235), .B1(n298), .B2(n256), .ZN(n296) );
  NAND2_X1 U303 ( .A1(n3), .A2(n341), .ZN(n298) );
  OAI22_X1 U304 ( .A1(n280), .A2(n235), .B1(n281), .B2(n256), .ZN(n279) );
  NOR3_X1 U305 ( .A1(n341), .A2(n280), .A3(n173), .ZN(n575) );
  NOR3_X1 U306 ( .A1(n341), .A2(n254), .A3(n173), .ZN(n563) );
  AOI21_X1 U307 ( .B1(n410), .B2(n16), .A(n511), .ZN(n505) );
  INV_X1 U308 ( .A(n507), .ZN(n511) );
  NOR3_X1 U309 ( .A1(n309), .A2(DATA2[3]), .A3(n310), .ZN(n308) );
  OAI21_X1 U310 ( .B1(n364), .B2(n353), .A(n535), .ZN(n492) );
  OAI21_X1 U311 ( .B1(n364), .B2(n339), .A(n174), .ZN(n149) );
  OAI21_X1 U312 ( .B1(n310), .B2(n20), .A(n507), .ZN(n231) );
  OAI21_X1 U313 ( .B1(n412), .B2(n353), .A(n658), .ZN(n307) );
  OAI21_X1 U314 ( .B1(n210), .B2(n20), .A(n632), .ZN(n302) );
  INV_X1 U315 ( .A(DATA2[4]), .ZN(n22) );
  NAND2_X1 U316 ( .A1(n12), .A2(n3), .ZN(n207) );
  OAI21_X1 U317 ( .B1(n364), .B2(n336), .A(n207), .ZN(n196) );
  NAND2_X1 U318 ( .A1(n145), .A2(n3), .ZN(n311) );
  AOI22_X1 U319 ( .A1(n229), .A2(n230), .B1(n231), .B2(n232), .ZN(n228) );
  NAND2_X1 U320 ( .A1(DATA2[3]), .A2(n3), .ZN(n174) );
  INV_X1 U321 ( .A(n3), .ZN(n233) );
  OAI211_X1 U322 ( .C1(n481), .C2(n22), .A(n482), .B(n483), .ZN(OUTSHFT[1]) );
  AOI21_X1 U323 ( .B1(n17), .B2(n488), .A(n489), .ZN(n482) );
  AOI22_X1 U324 ( .A1(n232), .A2(n491), .B1(n230), .B2(n492), .ZN(n481) );
  AOI221_X1 U325 ( .B1(n154), .B2(n484), .C1(n156), .C2(n485), .A(n486), .ZN(
        n483) );
  OAI211_X1 U326 ( .C1(n261), .C2(n22), .A(n262), .B(n263), .ZN(OUTSHFT[2]) );
  AOI21_X1 U327 ( .B1(n17), .B2(n269), .A(n270), .ZN(n262) );
  AOI22_X1 U328 ( .A1(n232), .A2(n272), .B1(n230), .B2(n273), .ZN(n261) );
  AOI221_X1 U329 ( .B1(n154), .B2(n264), .C1(n156), .C2(n265), .A(n266), .ZN(
        n263) );
  OAI21_X1 U330 ( .B1(n465), .B2(n466), .A(n467), .ZN(n464) );
  INV_X1 U331 ( .A(n204), .ZN(n465) );
  INV_X1 U332 ( .A(n627), .ZN(n361) );
  OAI221_X1 U333 ( .B1(n233), .B2(n579), .C1(n617), .C2(n8), .A(n335), .ZN(
        n627) );
  OAI21_X1 U334 ( .B1(n298), .B2(n309), .A(n311), .ZN(n306) );
  INV_X1 U335 ( .A(n703), .ZN(n432) );
  OAI221_X1 U336 ( .B1(n10), .B2(n28), .C1(n7), .C2(n29), .A(n704), .ZN(n703)
         );
  OAI21_X1 U337 ( .B1(n291), .B2(n219), .A(n248), .ZN(n290) );
  NAND2_X1 U338 ( .A1(n4), .A2(n3), .ZN(n234) );
  INV_X1 U339 ( .A(n669), .ZN(n402) );
  OAI221_X1 U340 ( .B1(n10), .B2(n33), .C1(n581), .C2(n34), .A(n671), .ZN(n669) );
  AOI22_X1 U341 ( .A1(DATA1[8]), .A2(n5), .B1(DATA1[7]), .B2(n4), .ZN(n671) );
  NAND4_X1 U342 ( .A1(n274), .A2(n248), .A3(n275), .A4(n276), .ZN(OUTSHFT[29])
         );
  OR2_X1 U343 ( .A1(n241), .A2(n284), .ZN(n274) );
  AOI22_X1 U344 ( .A1(n238), .A2(n282), .B1(n154), .B2(n283), .ZN(n275) );
  AOI221_X1 U345 ( .B1(n156), .B2(n277), .C1(n17), .C2(n278), .A(n279), .ZN(
        n276) );
  AOI22_X1 U346 ( .A1(n197), .A2(n150), .B1(n152), .B2(n198), .ZN(n191) );
  AOI221_X1 U347 ( .B1(n17), .B2(n193), .C1(n145), .C2(n194), .A(n195), .ZN(
        n192) );
  AOI22_X1 U348 ( .A1(n154), .A2(n199), .B1(n156), .B2(n200), .ZN(n190) );
  AOI22_X1 U349 ( .A1(n186), .A2(n150), .B1(n152), .B2(n187), .ZN(n180) );
  AOI221_X1 U350 ( .B1(n17), .B2(n182), .C1(n145), .C2(n183), .A(n184), .ZN(
        n181) );
  AOI22_X1 U351 ( .A1(n154), .A2(n188), .B1(n156), .B2(n189), .ZN(n179) );
  AOI22_X1 U352 ( .A1(n150), .A2(n151), .B1(n152), .B2(n153), .ZN(n141) );
  AOI221_X1 U353 ( .B1(n17), .B2(n144), .C1(n145), .C2(n146), .A(n147), .ZN(
        n142) );
  AOI22_X1 U354 ( .A1(n154), .A2(n155), .B1(n156), .B2(n157), .ZN(n140) );
  AOI22_X1 U355 ( .A1(n322), .A2(n150), .B1(n152), .B2(n326), .ZN(n679) );
  AOI221_X1 U356 ( .B1(n17), .B2(n325), .C1(n145), .C2(n328), .A(n681), .ZN(
        n680) );
  AOI22_X1 U357 ( .A1(n154), .A2(n327), .B1(n156), .B2(n321), .ZN(n678) );
  INV_X1 U358 ( .A(n584), .ZN(n6) );
  NAND2_X1 U359 ( .A1(n14), .A2(n359), .ZN(n354) );
  NAND2_X1 U360 ( .A1(n14), .A2(n436), .ZN(n683) );
  INV_X1 U361 ( .A(n479), .ZN(n387) );
  INV_X1 U362 ( .A(n460), .ZN(n360) );
  INV_X1 U363 ( .A(n510), .ZN(n411) );
  INV_X1 U364 ( .A(n225), .ZN(n230) );
  NAND2_X1 U365 ( .A1(n213), .A2(n214), .ZN(OUTSHFT[3]) );
  AOI221_X1 U366 ( .B1(n21), .B2(n222), .C1(n17), .C2(n223), .A(n224), .ZN(
        n213) );
  AOI221_X1 U367 ( .B1(n154), .B2(n215), .C1(n156), .C2(n216), .A(n217), .ZN(
        n214) );
  INV_X1 U368 ( .A(n228), .ZN(n222) );
  INV_X1 U369 ( .A(n386), .ZN(n297) );
  INV_X1 U370 ( .A(n440), .ZN(n523) );
  INV_X1 U371 ( .A(n502), .ZN(n396) );
  INV_X1 U372 ( .A(n478), .ZN(n373) );
  INV_X1 U373 ( .A(n405), .ZN(n555) );
  INV_X1 U374 ( .A(n472), .ZN(n372) );
  INV_X1 U375 ( .A(n509), .ZN(n397) );
  INV_X1 U376 ( .A(n381), .ZN(n634) );
  INV_X1 U377 ( .A(n451), .ZN(n338) );
  INV_X1 U378 ( .A(n346), .ZN(n449) );
  INV_X1 U379 ( .A(n376), .ZN(n470) );
  INV_X1 U380 ( .A(n459), .ZN(n340) );
  INV_X1 U381 ( .A(n525), .ZN(n423) );
  INV_X1 U382 ( .A(n684), .ZN(n325) );
  AOI221_X1 U383 ( .B1(n525), .B2(n15), .C1(n439), .C2(n14), .A(n685), .ZN(
        n684) );
  OAI22_X1 U384 ( .A1(n353), .A2(n517), .B1(n336), .B2(n422), .ZN(n685) );
  INV_X1 U385 ( .A(n576), .ZN(n281) );
  OAI21_X1 U386 ( .B1(n364), .B2(n341), .A(n298), .ZN(n576) );
  OR2_X1 U387 ( .A1(n241), .A2(n259), .ZN(n247) );
  AOI22_X1 U388 ( .A1(n260), .A2(n21), .B1(n22), .B2(n258), .ZN(n259) );
  OAI221_X1 U389 ( .B1(n615), .B2(n579), .C1(n617), .C2(n8), .A(n665), .ZN(
        n410) );
  AOI22_X1 U390 ( .A1(DATA1[28]), .A2(n5), .B1(DATA1[27]), .B2(n4), .ZN(n665)
         );
  OAI221_X1 U391 ( .B1(n10), .B2(n598), .C1(n592), .C2(n8), .A(n689), .ZN(n439) );
  AOI22_X1 U392 ( .A1(DATA1[25]), .A2(n5), .B1(DATA1[26]), .B2(n4), .ZN(n689)
         );
  OAI221_X1 U393 ( .B1(n10), .B2(n656), .C1(n9), .C2(n593), .A(n660), .ZN(n404) );
  AOI22_X1 U394 ( .A1(DATA1[20]), .A2(n5), .B1(DATA1[19]), .B2(n4), .ZN(n660)
         );
  OAI221_X1 U395 ( .B1(n579), .B2(n590), .C1(n8), .C2(n589), .A(n732), .ZN(
        n385) );
  AOI22_X1 U396 ( .A1(DATA1[25]), .A2(n5), .B1(DATA1[24]), .B2(n4), .ZN(n732)
         );
  OAI221_X1 U397 ( .B1(n10), .B2(n598), .C1(n581), .C2(n654), .A(n695), .ZN(
        n435) );
  OAI221_X1 U398 ( .B1(n10), .B2(n592), .C1(n9), .C2(n598), .A(n599), .ZN(n350) );
  OAI221_X1 U399 ( .B1(n579), .B2(n593), .C1(n592), .C2(n8), .A(n735), .ZN(
        n380) );
  AOI22_X1 U400 ( .A1(DATA1[21]), .A2(n584), .B1(DATA1[20]), .B2(n4), .ZN(n735) );
  OAI221_X1 U401 ( .B1(n579), .B2(n604), .C1(n581), .C2(n656), .A(n694), .ZN(
        n430) );
  AOI22_X1 U402 ( .A1(DATA1[19]), .A2(n5), .B1(DATA1[18]), .B2(n4), .ZN(n694)
         );
  OAI221_X1 U403 ( .B1(n579), .B2(n580), .C1(n9), .C2(n604), .A(n605), .ZN(
        n351) );
  OAI221_X1 U404 ( .B1(n10), .B2(n654), .C1(n8), .C2(n590), .A(n661), .ZN(n409) );
  AOI22_X1 U405 ( .A1(DATA1[24]), .A2(n5), .B1(DATA1[23]), .B2(n4), .ZN(n661)
         );
  OAI221_X1 U406 ( .B1(n10), .B2(n600), .C1(n615), .C2(n8), .A(n700), .ZN(n436) );
  AOI22_X1 U407 ( .A1(DATA1[27]), .A2(n5), .B1(DATA1[26]), .B2(n4), .ZN(n700)
         );
  OAI221_X1 U408 ( .B1(n10), .B2(n589), .C1(n9), .C2(n600), .A(n601), .ZN(n359) );
  AOI22_X1 U409 ( .A1(DATA1[26]), .A2(n584), .B1(DATA1[25]), .B2(n4), .ZN(n601) );
  OAI221_X1 U410 ( .B1(n617), .B2(n579), .C1(n233), .C2(n8), .A(n733), .ZN(
        n386) );
  AOI22_X1 U411 ( .A1(DATA1[29]), .A2(n5), .B1(DATA1[28]), .B2(n4), .ZN(n733)
         );
  OAI221_X1 U412 ( .B1(n10), .B2(n650), .C1(n8), .C2(n602), .A(n651), .ZN(n502) );
  AOI22_X1 U413 ( .A1(DATA1[18]), .A2(n5), .B1(DATA1[19]), .B2(n4), .ZN(n651)
         );
  OAI221_X1 U414 ( .B1(n10), .B2(n593), .C1(n7), .C2(n656), .A(n719), .ZN(n478) );
  AOI22_X1 U415 ( .A1(DATA1[23]), .A2(n5), .B1(DATA1[24]), .B2(n4), .ZN(n719)
         );
  OAI221_X1 U416 ( .B1(n10), .B2(n650), .C1(n8), .C2(n582), .A(n663), .ZN(n405) );
  AOI22_X1 U417 ( .A1(DATA1[16]), .A2(n5), .B1(DATA1[15]), .B2(n4), .ZN(n663)
         );
  OAI221_X1 U418 ( .B1(n10), .B2(n656), .C1(n8), .C2(n604), .A(n657), .ZN(n509) );
  OAI221_X1 U419 ( .B1(n579), .B2(n582), .C1(n7), .C2(n650), .A(n720), .ZN(
        n472) );
  AOI22_X1 U420 ( .A1(DATA1[19]), .A2(n5), .B1(DATA1[20]), .B2(n4), .ZN(n720)
         );
  OAI221_X1 U421 ( .B1(n579), .B2(n582), .C1(n8), .C2(n580), .A(n734), .ZN(
        n381) );
  OAI221_X1 U422 ( .B1(n10), .B2(n580), .C1(n9), .C2(n582), .A(n583), .ZN(n451) );
  AOI22_X1 U423 ( .A1(DATA1[20]), .A2(n584), .B1(DATA1[21]), .B2(n4), .ZN(n583) );
  OAI221_X1 U424 ( .B1(n8), .B2(n589), .C1(n6), .C2(n615), .A(n708), .ZN(n440)
         );
  AOI21_X1 U425 ( .B1(DATA1[28]), .B2(n11), .A(n682), .ZN(n708) );
  OAI221_X1 U426 ( .B1(n10), .B2(n38), .C1(n7), .C2(n37), .A(n716), .ZN(n376)
         );
  AOI22_X1 U427 ( .A1(DATA1[15]), .A2(n5), .B1(DATA1[16]), .B2(n4), .ZN(n716)
         );
  OAI221_X1 U428 ( .B1(n579), .B2(n2), .C1(n9), .C2(n38), .A(n588), .ZN(n346)
         );
  OAI221_X1 U429 ( .B1(n10), .B2(n592), .C1(n9), .C2(n593), .A(n594), .ZN(n459) );
  AOI22_X1 U430 ( .A1(DATA1[24]), .A2(n584), .B1(DATA1[25]), .B2(n4), .ZN(n594) );
  OAI221_X1 U431 ( .B1(n579), .B2(n604), .C1(n581), .C2(n580), .A(n690), .ZN(
        n525) );
  NAND2_X1 U432 ( .A1(n21), .A2(n493), .ZN(n173) );
  INV_X1 U433 ( .A(DATA1[29]), .ZN(n615) );
  INV_X1 U434 ( .A(DATA1[26]), .ZN(n590) );
  INV_X1 U435 ( .A(DATA1[25]), .ZN(n654) );
  OAI221_X1 U436 ( .B1(n10), .B2(n654), .C1(n8), .C2(n598), .A(n655), .ZN(n510) );
  AOI22_X1 U437 ( .A1(DATA1[26]), .A2(n5), .B1(DATA1[27]), .B2(n4), .ZN(n655)
         );
  OAI221_X1 U438 ( .B1(n10), .B2(n590), .C1(n7), .C2(n654), .A(n723), .ZN(n479) );
  AOI22_X1 U439 ( .A1(DATA1[27]), .A2(n5), .B1(DATA1[28]), .B2(n4), .ZN(n723)
         );
  OAI221_X1 U440 ( .B1(n579), .B2(n589), .C1(n9), .C2(n590), .A(n591), .ZN(
        n460) );
  AOI22_X1 U441 ( .A1(DATA1[28]), .A2(n584), .B1(DATA1[29]), .B2(n4), .ZN(n591) );
  INV_X1 U442 ( .A(DATA1[30]), .ZN(n617) );
  INV_X1 U443 ( .A(DATA1[18]), .ZN(n582) );
  INV_X1 U444 ( .A(DATA1[21]), .ZN(n656) );
  INV_X1 U445 ( .A(DATA1[28]), .ZN(n600) );
  INV_X1 U446 ( .A(DATA1[24]), .ZN(n598) );
  INV_X1 U447 ( .A(DATA1[20]), .ZN(n604) );
  INV_X1 U448 ( .A(DATA1[19]), .ZN(n580) );
  INV_X1 U449 ( .A(DATA1[27]), .ZN(n589) );
  INV_X1 U450 ( .A(DATA1[16]), .ZN(n602) );
  INV_X1 U451 ( .A(DATA1[23]), .ZN(n592) );
  AOI211_X1 U452 ( .C1(n225), .C2(n226), .A(n21), .B(n218), .ZN(n224) );
  AOI211_X1 U453 ( .C1(n225), .C2(n226), .A(n21), .B(n487), .ZN(n489) );
  AOI211_X1 U454 ( .C1(n225), .C2(n226), .A(n21), .B(n267), .ZN(n270) );
  OAI221_X1 U455 ( .B1(n709), .B2(n710), .C1(n370), .C2(n221), .A(n711), .ZN(
        OUTSHFT[0]) );
  NOR2_X1 U456 ( .A1(n692), .A2(n493), .ZN(n710) );
  AOI22_X1 U457 ( .A1(n21), .A2(n542), .B1(n543), .B2(n22), .ZN(n709) );
  AOI22_X1 U458 ( .A1(n154), .A2(n544), .B1(n17), .B2(n539), .ZN(n711) );
  OAI221_X1 U459 ( .B1(n233), .B2(n225), .C1(n234), .C2(n235), .A(n236), .ZN(
        OUTSHFT[31]) );
  AOI221_X1 U460 ( .B1(n156), .B2(n237), .C1(n238), .C2(n239), .A(n240), .ZN(
        n236) );
  AOI21_X1 U461 ( .B1(n241), .B2(n242), .A(n243), .ZN(n240) );
  AOI22_X1 U462 ( .A1(n21), .A2(n244), .B1(n245), .B2(n22), .ZN(n243) );
  NAND2_X1 U463 ( .A1(n692), .A2(n22), .ZN(n219) );
  NAND2_X1 U464 ( .A1(n493), .A2(n148), .ZN(n225) );
  NAND2_X1 U465 ( .A1(n493), .A2(n22), .ZN(n309) );
  NOR2_X1 U466 ( .A1(n242), .A2(n22), .ZN(n143) );
  NAND2_X1 U467 ( .A1(n299), .A2(n148), .ZN(n256) );
  NAND2_X1 U468 ( .A1(n292), .A2(n148), .ZN(n248) );
  NAND2_X1 U469 ( .A1(n692), .A2(n21), .ZN(n546) );
  INV_X1 U470 ( .A(DATA2[3]), .ZN(n20) );
  INV_X1 U471 ( .A(n226), .ZN(n232) );
  OAI211_X1 U472 ( .C1(n545), .C2(n546), .A(n547), .B(n548), .ZN(OUTSHFT[15])
         );
  INV_X1 U473 ( .A(n239), .ZN(n545) );
  AOI22_X1 U474 ( .A1(n237), .A2(n150), .B1(n314), .B2(n244), .ZN(n547) );
  AOI221_X1 U475 ( .B1(n292), .B2(n148), .C1(n17), .C2(n245), .A(n549), .ZN(
        n548) );
  INV_X1 U476 ( .A(n294), .ZN(n241) );
  INV_X1 U477 ( .A(n686), .ZN(n422) );
  OAI221_X1 U478 ( .B1(n10), .B2(n602), .C1(n581), .C2(n2), .A(n687), .ZN(n686) );
  AOI22_X1 U479 ( .A1(n208), .A2(n152), .B1(n209), .B2(n150), .ZN(n202) );
  AOI221_X1 U480 ( .B1(n17), .B2(n204), .C1(n145), .C2(n205), .A(n206), .ZN(
        n203) );
  AOI22_X1 U481 ( .A1(n154), .A2(n211), .B1(n156), .B2(n212), .ZN(n201) );
  AOI22_X1 U482 ( .A1(n175), .A2(n150), .B1(n152), .B2(n176), .ZN(n169) );
  AOI221_X1 U483 ( .B1(n17), .B2(n171), .C1(n145), .C2(n172), .A(n163), .ZN(
        n170) );
  AOI22_X1 U484 ( .A1(n154), .A2(n177), .B1(n156), .B2(n178), .ZN(n168) );
  AOI22_X1 U485 ( .A1(n164), .A2(n150), .B1(n152), .B2(n165), .ZN(n159) );
  AOI221_X1 U486 ( .B1(n17), .B2(n161), .C1(n145), .C2(n162), .A(n163), .ZN(
        n160) );
  AOI22_X1 U487 ( .A1(n154), .A2(n166), .B1(n156), .B2(n167), .ZN(n158) );
  AOI22_X1 U488 ( .A1(n317), .A2(n150), .B1(n152), .B2(n313), .ZN(n644) );
  AOI221_X1 U489 ( .B1(n17), .B2(n315), .C1(n646), .C2(n145), .A(n647), .ZN(
        n645) );
  AOI22_X1 U490 ( .A1(n154), .A2(n307), .B1(n156), .B2(n316), .ZN(n643) );
  AOI22_X1 U491 ( .A1(n277), .A2(n150), .B1(n152), .B2(n285), .ZN(n572) );
  AOI211_X1 U492 ( .C1(n17), .C2(n283), .A(n574), .B(n575), .ZN(n573) );
  AOI22_X1 U493 ( .A1(n154), .A2(n278), .B1(n156), .B2(n282), .ZN(n571) );
  AOI22_X1 U494 ( .A1(n251), .A2(n150), .B1(n152), .B2(n260), .ZN(n560) );
  AOI211_X1 U495 ( .C1(n17), .C2(n258), .A(n562), .B(n563), .ZN(n561) );
  AOI22_X1 U496 ( .A1(n154), .A2(n252), .B1(n156), .B2(n257), .ZN(n559) );
  INV_X1 U497 ( .A(n676), .ZN(n412) );
  OAI221_X1 U498 ( .B1(n8), .B2(n600), .C1(n6), .C2(n617), .A(n677), .ZN(n676)
         );
  AOI21_X1 U499 ( .B1(n11), .B2(DATA1[29]), .A(n648), .ZN(n677) );
  INV_X1 U500 ( .A(n721), .ZN(n388) );
  OAI221_X1 U501 ( .B1(n615), .B2(n8), .C1(n233), .C2(n6), .A(n722), .ZN(n721)
         );
  AOI21_X1 U502 ( .B1(n11), .B2(DATA1[30]), .A(n541), .ZN(n722) );
  NAND2_X1 U503 ( .A1(n286), .A2(n287), .ZN(OUTSHFT[28]) );
  AOI221_X1 U504 ( .B1(n17), .B2(n293), .C1(n294), .C2(n295), .A(n296), .ZN(
        n286) );
  AOI221_X1 U505 ( .B1(n154), .B2(n288), .C1(n156), .C2(n289), .A(n290), .ZN(
        n287) );
  INV_X1 U506 ( .A(n301), .ZN(n295) );
  AOI22_X1 U507 ( .A1(n238), .A2(n316), .B1(n156), .B2(n317), .ZN(n303) );
  AOI22_X1 U508 ( .A1(n312), .A2(n313), .B1(n314), .B2(n315), .ZN(n304) );
  AOI221_X1 U509 ( .B1(n306), .B2(n148), .C1(n17), .C2(n307), .A(n308), .ZN(
        n305) );
  CLKBUF_X1 U510 ( .A(DATA1[31]), .Z(n3) );
  AND3_X1 U511 ( .A1(n145), .A2(n148), .A3(n196), .ZN(n195) );
  AND3_X1 U512 ( .A1(n145), .A2(n148), .A3(n185), .ZN(n184) );
  AND3_X1 U513 ( .A1(n145), .A2(n148), .A3(n149), .ZN(n147) );
  AND3_X1 U514 ( .A1(n145), .A2(n148), .A3(n329), .ZN(n681) );
  NOR2_X1 U515 ( .A1(n39), .A2(FUNC[1]), .ZN(n493) );
  INV_X1 U516 ( .A(US), .ZN(n148) );
  NAND2_X1 U517 ( .A1(US), .A2(n493), .ZN(n226) );
  NOR3_X1 U518 ( .A1(n173), .A2(US), .A3(n174), .ZN(n163) );
  OAI211_X1 U519 ( .C1(US), .C2(n311), .A(n537), .B(n538), .ZN(OUTSHFT[16]) );
  AOI22_X1 U520 ( .A1(n156), .A2(n543), .B1(n17), .B2(n544), .ZN(n537) );
  AOI222_X1 U521 ( .A1(n539), .A2(n314), .B1(n540), .B2(n541), .C1(n542), .C2(
        n150), .ZN(n538) );
  INV_X1 U522 ( .A(n499), .ZN(n540) );
  OAI211_X1 U523 ( .C1(US), .C2(n526), .A(n527), .B(n528), .ZN(OUTSHFT[17]) );
  AOI21_X1 U524 ( .B1(n299), .B2(n492), .A(n292), .ZN(n526) );
  AOI22_X1 U525 ( .A1(n17), .A2(n484), .B1(n299), .B2(n491), .ZN(n527) );
  AOI221_X1 U526 ( .B1(n238), .B2(n485), .C1(n156), .C2(n490), .A(n529), .ZN(
        n528) );
  OAI211_X1 U527 ( .C1(US), .C2(n512), .A(n513), .B(n514), .ZN(OUTSHFT[18]) );
  AOI21_X1 U528 ( .B1(n299), .B2(n273), .A(n292), .ZN(n512) );
  AOI22_X1 U529 ( .A1(n17), .A2(n264), .B1(n299), .B2(n272), .ZN(n513) );
  AOI221_X1 U530 ( .B1(n238), .B2(n265), .C1(n156), .C2(n271), .A(n515), .ZN(
        n514) );
  OAI211_X1 U531 ( .C1(US), .C2(n494), .A(n495), .B(n496), .ZN(OUTSHFT[19]) );
  AOI21_X1 U532 ( .B1(n299), .B2(n229), .A(n292), .ZN(n494) );
  AOI22_X1 U533 ( .A1(n17), .A2(n215), .B1(n299), .B2(n231), .ZN(n495) );
  AOI221_X1 U534 ( .B1(n238), .B2(n216), .C1(n156), .C2(n227), .A(n497), .ZN(
        n496) );
  OAI211_X1 U535 ( .C1(US), .C2(n461), .A(n462), .B(n463), .ZN(OUTSHFT[20]) );
  AOI21_X1 U536 ( .B1(n299), .B2(n480), .A(n292), .ZN(n461) );
  AOI22_X1 U537 ( .A1(n17), .A2(n211), .B1(n299), .B2(n205), .ZN(n462) );
  AOI221_X1 U538 ( .B1(n238), .B2(n212), .C1(n156), .C2(n209), .A(n464), .ZN(
        n463) );
  OAI211_X1 U539 ( .C1(US), .C2(n443), .A(n444), .B(n445), .ZN(OUTSHFT[21]) );
  AOI21_X1 U540 ( .B1(n299), .B2(n196), .A(n292), .ZN(n443) );
  AOI22_X1 U541 ( .A1(n17), .A2(n199), .B1(n299), .B2(n194), .ZN(n444) );
  AOI221_X1 U542 ( .B1(n238), .B2(n200), .C1(n156), .C2(n197), .A(n446), .ZN(
        n445) );
  OAI211_X1 U543 ( .C1(US), .C2(n416), .A(n417), .B(n418), .ZN(OUTSHFT[22]) );
  AOI21_X1 U544 ( .B1(n299), .B2(n185), .A(n292), .ZN(n416) );
  AOI22_X1 U545 ( .A1(n17), .A2(n188), .B1(n299), .B2(n183), .ZN(n417) );
  AOI221_X1 U546 ( .B1(n238), .B2(n189), .C1(n156), .C2(n186), .A(n419), .ZN(
        n418) );
  OAI211_X1 U547 ( .C1(US), .C2(n365), .A(n391), .B(n392), .ZN(OUTSHFT[23]) );
  AOI22_X1 U549 ( .A1(n17), .A2(n177), .B1(n299), .B2(n172), .ZN(n391) );
  AOI221_X1 U550 ( .B1(n238), .B2(n178), .C1(n156), .C2(n175), .A(n393), .ZN(
        n392) );
  INV_X1 U552 ( .A(n394), .ZN(n393) );
  OAI211_X1 U553 ( .C1(US), .C2(n365), .A(n366), .B(n367), .ZN(OUTSHFT[24]) );
  AOI22_X1 U554 ( .A1(n17), .A2(n166), .B1(n299), .B2(n162), .ZN(n366) );
  AOI221_X1 U555 ( .B1(n238), .B2(n167), .C1(n156), .C2(n164), .A(n368), .ZN(
        n367) );
  INV_X1 U556 ( .A(n369), .ZN(n368) );
  OAI211_X1 U557 ( .C1(US), .C2(n330), .A(n331), .B(n332), .ZN(OUTSHFT[25]) );
  AOI21_X1 U558 ( .B1(n299), .B2(n149), .A(n292), .ZN(n330) );
  AOI22_X1 U559 ( .A1(n17), .A2(n155), .B1(n299), .B2(n146), .ZN(n331) );
  AOI221_X1 U560 ( .B1(n238), .B2(n157), .C1(n156), .C2(n151), .A(n333), .ZN(
        n332) );
  OAI211_X1 U561 ( .C1(US), .C2(n318), .A(n319), .B(n320), .ZN(OUTSHFT[26]) );
  AOI21_X1 U562 ( .B1(n299), .B2(n329), .A(n292), .ZN(n318) );
  AOI22_X1 U563 ( .A1(n17), .A2(n327), .B1(n299), .B2(n328), .ZN(n319) );
  AOI221_X1 U564 ( .B1(n238), .B2(n321), .C1(n156), .C2(n322), .A(n323), .ZN(
        n320) );
  NOR3_X1 U565 ( .A1(n173), .A2(US), .A3(n207), .ZN(n206) );
  NOR3_X1 U566 ( .A1(n173), .A2(US), .A3(n298), .ZN(n647) );
  NOR3_X1 U567 ( .A1(n173), .A2(US), .A3(n281), .ZN(n574) );
  NOR3_X1 U568 ( .A1(n173), .A2(US), .A3(n255), .ZN(n562) );
  NAND2_X1 U569 ( .A1(FUNC[1]), .A2(n39), .ZN(n242) );
  NOR2_X1 U570 ( .A1(FUNC[0]), .A2(FUNC[1]), .ZN(n294) );
  NAND4_X1 U571 ( .A1(n628), .A2(n629), .A3(n630), .A4(n631), .ZN(OUTSHFT[12])
         );
  OR3_X1 U572 ( .A1(n298), .A2(US), .A3(n173), .ZN(n629) );
  AOI22_X1 U573 ( .A1(n17), .A2(n288), .B1(n638), .B2(n145), .ZN(n628) );
  AOI22_X1 U574 ( .A1(n289), .A2(n150), .B1(n152), .B2(n302), .ZN(n631) );
  AND2_X1 U575 ( .A1(FUNC[1]), .A2(FUNC[0]), .ZN(n692) );
  NAND4_X1 U576 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(OUTSHFT[30])
         );
  INV_X1 U577 ( .A(DATA1[15]), .ZN(n2) );
  AOI22_X1 U578 ( .A1(DATA1[22]), .A2(n584), .B1(DATA1[21]), .B2(n4), .ZN(n599) );
  AOI22_X1 U579 ( .A1(DATA1[22]), .A2(n5), .B1(DATA1[23]), .B2(n4), .ZN(n657)
         );
  AOI22_X1 U580 ( .A1(DATA1[21]), .A2(n5), .B1(DATA1[22]), .B2(n4), .ZN(n690)
         );
  AOI22_X1 U581 ( .A1(DATA1[23]), .A2(n5), .B1(DATA1[22]), .B2(n4), .ZN(n695)
         );
  INV_X1 U582 ( .A(DATA1[22]), .ZN(n593) );
  AOI22_X1 U583 ( .A1(DATA1[16]), .A2(n584), .B1(DATA1[17]), .B2(n4), .ZN(n588) );
  AOI22_X1 U584 ( .A1(DATA1[18]), .A2(n5), .B1(DATA1[17]), .B2(n4), .ZN(n605)
         );
  AOI22_X1 U585 ( .A1(DATA1[17]), .A2(n5), .B1(DATA1[18]), .B2(n4), .ZN(n687)
         );
  AOI22_X1 U586 ( .A1(DATA1[17]), .A2(n5), .B1(DATA1[16]), .B2(n4), .ZN(n734)
         );
  INV_X1 U587 ( .A(DATA1[17]), .ZN(n650) );
  AOI22_X1 U588 ( .A1(DATA1[7]), .A2(n5), .B1(DATA1[6]), .B2(n4), .ZN(n701) );
  AOI22_X1 U589 ( .A1(DATA1[6]), .A2(n5), .B1(DATA1[7]), .B2(n4), .ZN(n675) );
  AOI22_X1 U590 ( .A1(n25), .A2(n584), .B1(DATA1[1]), .B2(n4), .ZN(n620) );
  AOI21_X1 U591 ( .B1(DATA1[1]), .B2(n11), .A(n648), .ZN(n666) );
  AOI22_X1 U592 ( .A1(DATA1[4]), .A2(n5), .B1(DATA1[5]), .B2(n4), .ZN(n624) );
  AOI22_X1 U593 ( .A1(DATA1[6]), .A2(n5), .B1(DATA1[5]), .B2(n4), .ZN(n609) );
  AOI22_X1 U594 ( .A1(DATA1[5]), .A2(n5), .B1(DATA1[6]), .B2(n4), .ZN(n705) );
  AOI22_X1 U595 ( .A1(DATA1[5]), .A2(n5), .B1(DATA1[4]), .B2(n4), .ZN(n727) );
  AOI22_X1 U596 ( .A1(DATA1[4]), .A2(n5), .B1(DATA1[3]), .B2(n4), .ZN(n668) );
  AOI22_X1 U597 ( .A1(n25), .A2(n5), .B1(DATA1[3]), .B2(n4), .ZN(n674) );
  AOI22_X1 U598 ( .A1(DATA1[3]), .A2(n5), .B1(n25), .B2(n4), .ZN(n704) );
  AOI22_X1 U599 ( .A1(DATA1[3]), .A2(n584), .B1(DATA1[4]), .B2(n4), .ZN(n715)
         );
  AOI22_X1 U600 ( .A1(n19), .A2(n410), .B1(DATA2[2]), .B2(n648), .ZN(n310) );
  OAI22_X1 U601 ( .A1(DATA2[2]), .A2(n476), .B1(n19), .B2(n370), .ZN(n468) );
  NAND2_X1 U602 ( .A1(DATA1[0]), .A2(n4), .ZN(n370) );
  AOI22_X1 U603 ( .A1(n4), .A2(DATA1[1]), .B1(n5), .B2(DATA1[0]), .ZN(n335) );
  NAND2_X1 U604 ( .A1(DATA2[1]), .A2(DATA2[0]), .ZN(n581) );
  NAND2_X1 U605 ( .A1(DATA2[1]), .A2(n18), .ZN(n579) );
  NOR2_X1 U606 ( .A1(n18), .A2(DATA2[1]), .ZN(n584) );
  AOI21_X1 U607 ( .B1(n3), .B2(DATA2[1]), .A(n577), .ZN(n364) );
  INV_X1 U608 ( .A(n579), .ZN(n11) );
  INV_X1 U609 ( .A(DATA2[0]), .ZN(n18) );
  INV_X1 U610 ( .A(DATA2[2]), .ZN(n19) );
  INV_X1 U611 ( .A(n22), .ZN(n21) );
  INV_X1 U612 ( .A(DATA1[0]), .ZN(n23) );
  INV_X1 U613 ( .A(DATA1[1]), .ZN(n24) );
  INV_X1 U614 ( .A(n26), .ZN(n25) );
  INV_X1 U615 ( .A(DATA1[2]), .ZN(n26) );
  INV_X1 U616 ( .A(DATA1[3]), .ZN(n27) );
  INV_X1 U617 ( .A(DATA1[4]), .ZN(n28) );
  INV_X1 U618 ( .A(DATA1[5]), .ZN(n29) );
  INV_X1 U631 ( .A(DATA1[6]), .ZN(n30) );
  INV_X1 U632 ( .A(DATA1[7]), .ZN(n31) );
  INV_X1 U633 ( .A(DATA1[8]), .ZN(n32) );
  INV_X1 U634 ( .A(DATA1[9]), .ZN(n33) );
  INV_X1 U635 ( .A(DATA1[10]), .ZN(n34) );
  INV_X1 U636 ( .A(DATA1[11]), .ZN(n35) );
  INV_X1 U637 ( .A(DATA1[12]), .ZN(n36) );
  INV_X1 U638 ( .A(DATA1[13]), .ZN(n37) );
  INV_X1 U639 ( .A(DATA1[14]), .ZN(n38) );
  INV_X1 U640 ( .A(FUNC[0]), .ZN(n39) );
endmodule


module BOOTHMUL_NB32_0 ( A, B, C );
  input [15:0] A;
  input [15:0] B;
  output [31:0] C;
  wire   \Term[7][31] , \Term[7][30] , \Term[7][29] , \Term[7][28] ,
         \Term[7][27] , \Term[7][26] , \Term[7][25] , \Term[7][24] ,
         \Term[7][23] , \Term[7][22] , \Term[7][21] , \Term[7][20] ,
         \Term[7][19] , \Term[7][18] , \Term[7][17] , \Term[7][16] ,
         \Term[7][15] , \Term[7][14] , \Term[7][13] , \Term[7][12] ,
         \Term[7][11] , \Term[7][10] , \Term[7][9] , \Term[7][8] ,
         \Term[7][7] , \Term[7][6] , \Term[7][5] , \Term[7][4] , \Term[7][3] ,
         \Term[7][2] , \Term[7][1] , \Term[7][0] , \Term[6][31] ,
         \Term[6][30] , \Term[6][29] , \Term[6][28] , \Term[6][27] ,
         \Term[6][26] , \Term[6][25] , \Term[6][24] , \Term[6][23] ,
         \Term[6][22] , \Term[6][21] , \Term[6][20] , \Term[6][19] ,
         \Term[6][18] , \Term[6][17] , \Term[6][16] , \Term[6][15] ,
         \Term[6][14] , \Term[6][13] , \Term[6][12] , \Term[6][11] ,
         \Term[6][10] , \Term[6][9] , \Term[6][8] , \Term[6][7] , \Term[6][6] ,
         \Term[6][5] , \Term[6][4] , \Term[6][3] , \Term[6][2] , \Term[6][1] ,
         \Term[6][0] , \Term[5][31] , \Term[5][30] , \Term[5][29] ,
         \Term[5][28] , \Term[5][27] , \Term[5][26] , \Term[5][25] ,
         \Term[5][24] , \Term[5][23] , \Term[5][22] , \Term[5][21] ,
         \Term[5][20] , \Term[5][19] , \Term[5][18] , \Term[5][17] ,
         \Term[5][16] , \Term[5][15] , \Term[5][14] , \Term[5][13] ,
         \Term[5][12] , \Term[5][11] , \Term[5][10] , \Term[5][9] ,
         \Term[5][8] , \Term[5][7] , \Term[5][6] , \Term[5][5] , \Term[5][4] ,
         \Term[5][3] , \Term[5][2] , \Term[5][1] , \Term[5][0] , \Term[4][31] ,
         \Term[4][30] , \Term[4][29] , \Term[4][28] , \Term[4][27] ,
         \Term[4][26] , \Term[4][25] , \Term[4][24] , \Term[4][23] ,
         \Term[4][22] , \Term[4][21] , \Term[4][20] , \Term[4][19] ,
         \Term[4][18] , \Term[4][17] , \Term[4][16] , \Term[4][15] ,
         \Term[4][14] , \Term[4][13] , \Term[4][12] , \Term[4][11] ,
         \Term[4][10] , \Term[4][9] , \Term[4][8] , \Term[4][7] , \Term[4][6] ,
         \Term[4][5] , \Term[4][4] , \Term[4][3] , \Term[4][2] , \Term[4][1] ,
         \Term[4][0] , \Term[3][31] , \Term[3][30] , \Term[3][29] ,
         \Term[3][28] , \Term[3][27] , \Term[3][26] , \Term[3][25] ,
         \Term[3][24] , \Term[3][23] , \Term[3][22] , \Term[3][21] ,
         \Term[3][20] , \Term[3][19] , \Term[3][18] , \Term[3][17] ,
         \Term[3][16] , \Term[3][15] , \Term[3][14] , \Term[3][13] ,
         \Term[3][12] , \Term[3][11] , \Term[3][10] , \Term[3][9] ,
         \Term[3][8] , \Term[3][7] , \Term[3][6] , \Term[3][5] , \Term[3][4] ,
         \Term[3][3] , \Term[3][2] , \Term[3][1] , \Term[3][0] , \Term[2][31] ,
         \Term[2][30] , \Term[2][29] , \Term[2][28] , \Term[2][27] ,
         \Term[2][26] , \Term[2][25] , \Term[2][24] , \Term[2][23] ,
         \Term[2][22] , \Term[2][21] , \Term[2][20] , \Term[2][19] ,
         \Term[2][18] , \Term[2][17] , \Term[2][16] , \Term[2][15] ,
         \Term[2][14] , \Term[2][13] , \Term[2][12] , \Term[2][11] ,
         \Term[2][10] , \Term[2][9] , \Term[2][8] , \Term[2][7] , \Term[2][6] ,
         \Term[2][5] , \Term[2][4] , \Term[2][3] , \Term[2][2] , \Term[2][1] ,
         \Term[2][0] , \Term[1][31] , \Term[1][30] , \Term[1][29] ,
         \Term[1][28] , \Term[1][27] , \Term[1][26] , \Term[1][25] ,
         \Term[1][24] , \Term[1][23] , \Term[1][22] , \Term[1][21] ,
         \Term[1][20] , \Term[1][19] , \Term[1][18] , \Term[1][17] ,
         \Term[1][16] , \Term[1][15] , \Term[1][14] , \Term[1][13] ,
         \Term[1][12] , \Term[1][11] , \Term[1][10] , \Term[1][9] ,
         \Term[1][8] , \Term[1][7] , \Term[1][6] , \Term[1][5] , \Term[1][4] ,
         \Term[1][3] , \Term[1][2] , \Term[1][1] , \Term[1][0] , \Term[0][31] ,
         \Term[0][30] , \Term[0][29] , \Term[0][28] , \Term[0][27] ,
         \Term[0][26] , \Term[0][25] , \Term[0][24] , \Term[0][23] ,
         \Term[0][22] , \Term[0][21] , \Term[0][20] , \Term[0][19] ,
         \Term[0][18] , \Term[0][17] , \Term[0][16] , \Term[0][15] ,
         \Term[0][14] , \Term[0][13] , \Term[0][12] , \Term[0][11] ,
         \Term[0][10] , \Term[0][9] , \Term[0][8] , \Term[0][7] , \Term[0][6] ,
         \Term[0][5] , \Term[0][4] , \Term[0][3] , \Term[0][2] , \Term[0][1] ,
         \Term[0][0] , \Res[6][31] , \Res[6][30] , \Res[6][29] , \Res[6][28] ,
         \Res[6][27] , \Res[6][26] , \Res[6][25] , \Res[6][24] , \Res[6][23] ,
         \Res[6][22] , \Res[6][21] , \Res[6][20] , \Res[6][19] , \Res[6][18] ,
         \Res[6][17] , \Res[6][16] , \Res[6][15] , \Res[6][14] , \Res[6][13] ,
         \Res[6][12] , \Res[6][11] , \Res[6][10] , \Res[6][9] , \Res[6][8] ,
         \Res[6][7] , \Res[6][6] , \Res[6][5] , \Res[6][4] , \Res[6][3] ,
         \Res[6][2] , \Res[6][1] , \Res[6][0] , \Res[5][31] , \Res[5][30] ,
         \Res[5][29] , \Res[5][28] , \Res[5][27] , \Res[5][26] , \Res[5][25] ,
         \Res[5][24] , \Res[5][23] , \Res[5][22] , \Res[5][21] , \Res[5][20] ,
         \Res[5][19] , \Res[5][18] , \Res[5][17] , \Res[5][16] , \Res[5][15] ,
         \Res[5][14] , \Res[5][13] , \Res[5][12] , \Res[5][11] , \Res[5][10] ,
         \Res[5][9] , \Res[5][8] , \Res[5][7] , \Res[5][6] , \Res[5][5] ,
         \Res[5][4] , \Res[5][3] , \Res[5][2] , \Res[5][1] , \Res[5][0] ,
         \Res[4][31] , \Res[4][30] , \Res[4][29] , \Res[4][28] , \Res[4][27] ,
         \Res[4][26] , \Res[4][25] , \Res[4][24] , \Res[4][23] , \Res[4][22] ,
         \Res[4][21] , \Res[4][20] , \Res[4][19] , \Res[4][18] , \Res[4][17] ,
         \Res[4][16] , \Res[4][15] , \Res[4][14] , \Res[4][13] , \Res[4][12] ,
         \Res[4][11] , \Res[4][10] , \Res[4][9] , \Res[4][8] , \Res[4][7] ,
         \Res[4][6] , \Res[4][5] , \Res[4][4] , \Res[4][3] , \Res[4][2] ,
         \Res[4][1] , \Res[4][0] , \Res[3][31] , \Res[3][30] , \Res[3][29] ,
         \Res[3][28] , \Res[3][27] , \Res[3][26] , \Res[3][25] , \Res[3][24] ,
         \Res[3][23] , \Res[3][22] , \Res[3][21] , \Res[3][20] , \Res[3][19] ,
         \Res[3][18] , \Res[3][17] , \Res[3][16] , \Res[3][15] , \Res[3][14] ,
         \Res[3][13] , \Res[3][12] , \Res[3][11] , \Res[3][10] , \Res[3][9] ,
         \Res[3][8] , \Res[3][7] , \Res[3][6] , \Res[3][5] , \Res[3][4] ,
         \Res[3][3] , \Res[3][2] , \Res[3][1] , \Res[3][0] , \Res[2][31] ,
         \Res[2][30] , \Res[2][29] , \Res[2][28] , \Res[2][27] , \Res[2][26] ,
         \Res[2][25] , \Res[2][24] , \Res[2][23] , \Res[2][22] , \Res[2][21] ,
         \Res[2][20] , \Res[2][19] , \Res[2][18] , \Res[2][17] , \Res[2][16] ,
         \Res[2][15] , \Res[2][14] , \Res[2][13] , \Res[2][12] , \Res[2][11] ,
         \Res[2][10] , \Res[2][9] , \Res[2][8] , \Res[2][7] , \Res[2][6] ,
         \Res[2][5] , \Res[2][4] , \Res[2][3] , \Res[2][2] , \Res[2][1] ,
         \Res[2][0] , \Res[1][31] , \Res[1][30] , \Res[1][29] , \Res[1][28] ,
         \Res[1][27] , \Res[1][26] , \Res[1][25] , \Res[1][24] , \Res[1][23] ,
         \Res[1][22] , \Res[1][21] , \Res[1][20] , \Res[1][19] , \Res[1][18] ,
         \Res[1][17] , \Res[1][16] , \Res[1][15] , \Res[1][14] , \Res[1][13] ,
         \Res[1][12] , \Res[1][11] , \Res[1][10] , \Res[1][9] , \Res[1][8] ,
         \Res[1][7] , \Res[1][6] , \Res[1][5] , \Res[1][4] , \Res[1][3] ,
         \Res[1][2] , \Res[1][1] , \Res[1][0] , \Res[0][31] , \Res[0][30] ,
         \Res[0][29] , \Res[0][28] , \Res[0][27] , \Res[0][26] , \Res[0][25] ,
         \Res[0][24] , \Res[0][23] , \Res[0][22] , \Res[0][21] , \Res[0][20] ,
         \Res[0][19] , \Res[0][18] , \Res[0][17] , \Res[0][16] , \Res[0][15] ,
         \Res[0][14] , \Res[0][13] , \Res[0][12] , \Res[0][11] , \Res[0][10] ,
         \Res[0][9] , \Res[0][8] , \Res[0][7] , \Res[0][6] , \Res[0][5] ,
         \Res[0][4] , \Res[0][3] , \Res[0][2] , \Res[0][1] , \Res[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [7:0] OP;

  CLKBUF_X1 U2 ( .A(A[8]), .Z(n8) );
  CLKBUF_X1 U3 ( .A(A[12]), .Z(n12) );
  CLKBUF_X1 U4 ( .A(A[11]), .Z(n11) );
  CLKBUF_X1 U5 ( .A(A[9]), .Z(n9) );
  CLKBUF_X1 U6 ( .A(A[10]), .Z(n10) );
  CLKBUF_X1 U7 ( .A(A[13]), .Z(n13) );
  CLKBUF_X1 U8 ( .A(A[14]), .Z(n14) );
  CLKBUF_X1 U9 ( .A(A[7]), .Z(n7) );
  CLKBUF_X1 U10 ( .A(A[4]), .Z(n4) );
  CLKBUF_X1 U11 ( .A(A[5]), .Z(n5) );
  CLKBUF_X1 U12 ( .A(A[6]), .Z(n6) );
  CLKBUF_X1 U13 ( .A(A[2]), .Z(n2) );
  CLKBUF_X1 U14 ( .A(A[1]), .Z(n1) );
  CLKBUF_X1 U15 ( .A(A[3]), .Z(n3) );
  MUX_SHIFT_NB16_N_sh0_0 mux_map_0 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel({B[1:0], 1'b0}), .AS(
        OP[0]), .B({\Term[0][31] , \Term[0][30] , \Term[0][29] , \Term[0][28] , 
        \Term[0][27] , \Term[0][26] , \Term[0][25] , \Term[0][24] , 
        \Term[0][23] , \Term[0][22] , \Term[0][21] , \Term[0][20] , 
        \Term[0][19] , \Term[0][18] , \Term[0][17] , \Term[0][16] , 
        \Term[0][15] , \Term[0][14] , \Term[0][13] , \Term[0][12] , 
        \Term[0][11] , \Term[0][10] , \Term[0][9] , \Term[0][8] , \Term[0][7] , 
        \Term[0][6] , \Term[0][5] , \Term[0][4] , \Term[0][3] , \Term[0][2] , 
        \Term[0][1] , \Term[0][0] }) );
  MUX_SHIFT_NB16_N_sh2_0 mux_map_1 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel(B[3:1]), .AS(OP[1]), .B({
        \Term[1][31] , \Term[1][30] , \Term[1][29] , \Term[1][28] , 
        \Term[1][27] , \Term[1][26] , \Term[1][25] , \Term[1][24] , 
        \Term[1][23] , \Term[1][22] , \Term[1][21] , \Term[1][20] , 
        \Term[1][19] , \Term[1][18] , \Term[1][17] , \Term[1][16] , 
        \Term[1][15] , \Term[1][14] , \Term[1][13] , \Term[1][12] , 
        \Term[1][11] , \Term[1][10] , \Term[1][9] , \Term[1][8] , \Term[1][7] , 
        \Term[1][6] , \Term[1][5] , \Term[1][4] , \Term[1][3] , \Term[1][2] , 
        \Term[1][1] , \Term[1][0] }) );
  MUX_SHIFT_NB16_N_sh4_0 mux_map_2 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel(B[5:3]), .AS(OP[2]), .B({
        \Term[2][31] , \Term[2][30] , \Term[2][29] , \Term[2][28] , 
        \Term[2][27] , \Term[2][26] , \Term[2][25] , \Term[2][24] , 
        \Term[2][23] , \Term[2][22] , \Term[2][21] , \Term[2][20] , 
        \Term[2][19] , \Term[2][18] , \Term[2][17] , \Term[2][16] , 
        \Term[2][15] , \Term[2][14] , \Term[2][13] , \Term[2][12] , 
        \Term[2][11] , \Term[2][10] , \Term[2][9] , \Term[2][8] , \Term[2][7] , 
        \Term[2][6] , \Term[2][5] , \Term[2][4] , \Term[2][3] , \Term[2][2] , 
        \Term[2][1] , \Term[2][0] }) );
  MUX_SHIFT_NB16_N_sh6_0 mux_map_3 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel(B[7:5]), .AS(OP[3]), .B({
        \Term[3][31] , \Term[3][30] , \Term[3][29] , \Term[3][28] , 
        \Term[3][27] , \Term[3][26] , \Term[3][25] , \Term[3][24] , 
        \Term[3][23] , \Term[3][22] , \Term[3][21] , \Term[3][20] , 
        \Term[3][19] , \Term[3][18] , \Term[3][17] , \Term[3][16] , 
        \Term[3][15] , \Term[3][14] , \Term[3][13] , \Term[3][12] , 
        \Term[3][11] , \Term[3][10] , \Term[3][9] , \Term[3][8] , \Term[3][7] , 
        \Term[3][6] , \Term[3][5] , \Term[3][4] , \Term[3][3] , \Term[3][2] , 
        \Term[3][1] , \Term[3][0] }) );
  MUX_SHIFT_NB16_N_sh8_0 mux_map_4 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel(B[9:7]), .AS(OP[4]), .B({
        \Term[4][31] , \Term[4][30] , \Term[4][29] , \Term[4][28] , 
        \Term[4][27] , \Term[4][26] , \Term[4][25] , \Term[4][24] , 
        \Term[4][23] , \Term[4][22] , \Term[4][21] , \Term[4][20] , 
        \Term[4][19] , \Term[4][18] , \Term[4][17] , \Term[4][16] , 
        \Term[4][15] , \Term[4][14] , \Term[4][13] , \Term[4][12] , 
        \Term[4][11] , \Term[4][10] , \Term[4][9] , \Term[4][8] , \Term[4][7] , 
        \Term[4][6] , \Term[4][5] , \Term[4][4] , \Term[4][3] , \Term[4][2] , 
        \Term[4][1] , \Term[4][0] }) );
  MUX_SHIFT_NB16_N_sh10_0 mux_map_5 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel(B[11:9]), .AS(OP[5]), .B(
        {\Term[5][31] , \Term[5][30] , \Term[5][29] , \Term[5][28] , 
        \Term[5][27] , \Term[5][26] , \Term[5][25] , \Term[5][24] , 
        \Term[5][23] , \Term[5][22] , \Term[5][21] , \Term[5][20] , 
        \Term[5][19] , \Term[5][18] , \Term[5][17] , \Term[5][16] , 
        \Term[5][15] , \Term[5][14] , \Term[5][13] , \Term[5][12] , 
        \Term[5][11] , \Term[5][10] , \Term[5][9] , \Term[5][8] , \Term[5][7] , 
        \Term[5][6] , \Term[5][5] , \Term[5][4] , \Term[5][3] , \Term[5][2] , 
        \Term[5][1] , \Term[5][0] }) );
  MUX_SHIFT_NB16_N_sh12_0 mux_map_6 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel(B[13:11]), .AS(OP[6]), 
        .B({\Term[6][31] , \Term[6][30] , \Term[6][29] , \Term[6][28] , 
        \Term[6][27] , \Term[6][26] , \Term[6][25] , \Term[6][24] , 
        \Term[6][23] , \Term[6][22] , \Term[6][21] , \Term[6][20] , 
        \Term[6][19] , \Term[6][18] , \Term[6][17] , \Term[6][16] , 
        \Term[6][15] , \Term[6][14] , \Term[6][13] , \Term[6][12] , 
        \Term[6][11] , \Term[6][10] , \Term[6][9] , \Term[6][8] , \Term[6][7] , 
        \Term[6][6] , \Term[6][5] , \Term[6][4] , \Term[6][3] , \Term[6][2] , 
        \Term[6][1] , \Term[6][0] }) );
  MUX_SHIFT_NB16_N_sh14_0 mux_map_7 ( .A({A[15], n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1, A[0]}), .sel(B[15:13]), .AS(OP[7]), 
        .B({\Term[7][31] , \Term[7][30] , \Term[7][29] , \Term[7][28] , 
        \Term[7][27] , \Term[7][26] , \Term[7][25] , \Term[7][24] , 
        \Term[7][23] , \Term[7][22] , \Term[7][21] , \Term[7][20] , 
        \Term[7][19] , \Term[7][18] , \Term[7][17] , \Term[7][16] , 
        \Term[7][15] , \Term[7][14] , \Term[7][13] , \Term[7][12] , 
        \Term[7][11] , \Term[7][10] , \Term[7][9] , \Term[7][8] , \Term[7][7] , 
        \Term[7][6] , \Term[7][5] , \Term[7][4] , \Term[7][3] , \Term[7][2] , 
        \Term[7][1] , \Term[7][0] }) );
  p4addgen_NB32_CW4_7 adder_0 ( .A({\Term[0][31] , \Term[0][30] , 
        \Term[0][29] , \Term[0][28] , \Term[0][27] , \Term[0][26] , 
        \Term[0][25] , \Term[0][24] , \Term[0][23] , \Term[0][22] , 
        \Term[0][21] , \Term[0][20] , \Term[0][19] , \Term[0][18] , 
        \Term[0][17] , \Term[0][16] , \Term[0][15] , \Term[0][14] , 
        \Term[0][13] , \Term[0][12] , \Term[0][11] , \Term[0][10] , 
        \Term[0][9] , \Term[0][8] , \Term[0][7] , \Term[0][6] , \Term[0][5] , 
        \Term[0][4] , \Term[0][3] , \Term[0][2] , \Term[0][1] , \Term[0][0] }), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Ci(OP[0]), 
        .S({\Res[0][31] , \Res[0][30] , \Res[0][29] , \Res[0][28] , 
        \Res[0][27] , \Res[0][26] , \Res[0][25] , \Res[0][24] , \Res[0][23] , 
        \Res[0][22] , \Res[0][21] , \Res[0][20] , \Res[0][19] , \Res[0][18] , 
        \Res[0][17] , \Res[0][16] , \Res[0][15] , \Res[0][14] , \Res[0][13] , 
        \Res[0][12] , \Res[0][11] , \Res[0][10] , \Res[0][9] , \Res[0][8] , 
        \Res[0][7] , \Res[0][6] , \Res[0][5] , \Res[0][4] , \Res[0][3] , 
        \Res[0][2] , \Res[0][1] , \Res[0][0] }) );
  p4addgen_NB32_CW4_6 add_map_1 ( .A({\Term[1][31] , \Term[1][30] , 
        \Term[1][29] , \Term[1][28] , \Term[1][27] , \Term[1][26] , 
        \Term[1][25] , \Term[1][24] , \Term[1][23] , \Term[1][22] , 
        \Term[1][21] , \Term[1][20] , \Term[1][19] , \Term[1][18] , 
        \Term[1][17] , \Term[1][16] , \Term[1][15] , \Term[1][14] , 
        \Term[1][13] , \Term[1][12] , \Term[1][11] , \Term[1][10] , 
        \Term[1][9] , \Term[1][8] , \Term[1][7] , \Term[1][6] , \Term[1][5] , 
        \Term[1][4] , \Term[1][3] , \Term[1][2] , \Term[1][1] , \Term[1][0] }), 
        .B({\Res[0][31] , \Res[0][30] , \Res[0][29] , \Res[0][28] , 
        \Res[0][27] , \Res[0][26] , \Res[0][25] , \Res[0][24] , \Res[0][23] , 
        \Res[0][22] , \Res[0][21] , \Res[0][20] , \Res[0][19] , \Res[0][18] , 
        \Res[0][17] , \Res[0][16] , \Res[0][15] , \Res[0][14] , \Res[0][13] , 
        \Res[0][12] , \Res[0][11] , \Res[0][10] , \Res[0][9] , \Res[0][8] , 
        \Res[0][7] , \Res[0][6] , \Res[0][5] , \Res[0][4] , \Res[0][3] , 
        \Res[0][2] , \Res[0][1] , \Res[0][0] }), .Ci(OP[1]), .S({\Res[1][31] , 
        \Res[1][30] , \Res[1][29] , \Res[1][28] , \Res[1][27] , \Res[1][26] , 
        \Res[1][25] , \Res[1][24] , \Res[1][23] , \Res[1][22] , \Res[1][21] , 
        \Res[1][20] , \Res[1][19] , \Res[1][18] , \Res[1][17] , \Res[1][16] , 
        \Res[1][15] , \Res[1][14] , \Res[1][13] , \Res[1][12] , \Res[1][11] , 
        \Res[1][10] , \Res[1][9] , \Res[1][8] , \Res[1][7] , \Res[1][6] , 
        \Res[1][5] , \Res[1][4] , \Res[1][3] , \Res[1][2] , \Res[1][1] , 
        \Res[1][0] }) );
  p4addgen_NB32_CW4_5 add_map_2 ( .A({\Term[2][31] , \Term[2][30] , 
        \Term[2][29] , \Term[2][28] , \Term[2][27] , \Term[2][26] , 
        \Term[2][25] , \Term[2][24] , \Term[2][23] , \Term[2][22] , 
        \Term[2][21] , \Term[2][20] , \Term[2][19] , \Term[2][18] , 
        \Term[2][17] , \Term[2][16] , \Term[2][15] , \Term[2][14] , 
        \Term[2][13] , \Term[2][12] , \Term[2][11] , \Term[2][10] , 
        \Term[2][9] , \Term[2][8] , \Term[2][7] , \Term[2][6] , \Term[2][5] , 
        \Term[2][4] , \Term[2][3] , \Term[2][2] , \Term[2][1] , \Term[2][0] }), 
        .B({\Res[1][31] , \Res[1][30] , \Res[1][29] , \Res[1][28] , 
        \Res[1][27] , \Res[1][26] , \Res[1][25] , \Res[1][24] , \Res[1][23] , 
        \Res[1][22] , \Res[1][21] , \Res[1][20] , \Res[1][19] , \Res[1][18] , 
        \Res[1][17] , \Res[1][16] , \Res[1][15] , \Res[1][14] , \Res[1][13] , 
        \Res[1][12] , \Res[1][11] , \Res[1][10] , \Res[1][9] , \Res[1][8] , 
        \Res[1][7] , \Res[1][6] , \Res[1][5] , \Res[1][4] , \Res[1][3] , 
        \Res[1][2] , \Res[1][1] , \Res[1][0] }), .Ci(OP[2]), .S({\Res[2][31] , 
        \Res[2][30] , \Res[2][29] , \Res[2][28] , \Res[2][27] , \Res[2][26] , 
        \Res[2][25] , \Res[2][24] , \Res[2][23] , \Res[2][22] , \Res[2][21] , 
        \Res[2][20] , \Res[2][19] , \Res[2][18] , \Res[2][17] , \Res[2][16] , 
        \Res[2][15] , \Res[2][14] , \Res[2][13] , \Res[2][12] , \Res[2][11] , 
        \Res[2][10] , \Res[2][9] , \Res[2][8] , \Res[2][7] , \Res[2][6] , 
        \Res[2][5] , \Res[2][4] , \Res[2][3] , \Res[2][2] , \Res[2][1] , 
        \Res[2][0] }) );
  p4addgen_NB32_CW4_4 add_map_3 ( .A({\Term[3][31] , \Term[3][30] , 
        \Term[3][29] , \Term[3][28] , \Term[3][27] , \Term[3][26] , 
        \Term[3][25] , \Term[3][24] , \Term[3][23] , \Term[3][22] , 
        \Term[3][21] , \Term[3][20] , \Term[3][19] , \Term[3][18] , 
        \Term[3][17] , \Term[3][16] , \Term[3][15] , \Term[3][14] , 
        \Term[3][13] , \Term[3][12] , \Term[3][11] , \Term[3][10] , 
        \Term[3][9] , \Term[3][8] , \Term[3][7] , \Term[3][6] , \Term[3][5] , 
        \Term[3][4] , \Term[3][3] , \Term[3][2] , \Term[3][1] , \Term[3][0] }), 
        .B({\Res[2][31] , \Res[2][30] , \Res[2][29] , \Res[2][28] , 
        \Res[2][27] , \Res[2][26] , \Res[2][25] , \Res[2][24] , \Res[2][23] , 
        \Res[2][22] , \Res[2][21] , \Res[2][20] , \Res[2][19] , \Res[2][18] , 
        \Res[2][17] , \Res[2][16] , \Res[2][15] , \Res[2][14] , \Res[2][13] , 
        \Res[2][12] , \Res[2][11] , \Res[2][10] , \Res[2][9] , \Res[2][8] , 
        \Res[2][7] , \Res[2][6] , \Res[2][5] , \Res[2][4] , \Res[2][3] , 
        \Res[2][2] , \Res[2][1] , \Res[2][0] }), .Ci(OP[3]), .S({\Res[3][31] , 
        \Res[3][30] , \Res[3][29] , \Res[3][28] , \Res[3][27] , \Res[3][26] , 
        \Res[3][25] , \Res[3][24] , \Res[3][23] , \Res[3][22] , \Res[3][21] , 
        \Res[3][20] , \Res[3][19] , \Res[3][18] , \Res[3][17] , \Res[3][16] , 
        \Res[3][15] , \Res[3][14] , \Res[3][13] , \Res[3][12] , \Res[3][11] , 
        \Res[3][10] , \Res[3][9] , \Res[3][8] , \Res[3][7] , \Res[3][6] , 
        \Res[3][5] , \Res[3][4] , \Res[3][3] , \Res[3][2] , \Res[3][1] , 
        \Res[3][0] }) );
  p4addgen_NB32_CW4_3 add_map_4 ( .A({\Term[4][31] , \Term[4][30] , 
        \Term[4][29] , \Term[4][28] , \Term[4][27] , \Term[4][26] , 
        \Term[4][25] , \Term[4][24] , \Term[4][23] , \Term[4][22] , 
        \Term[4][21] , \Term[4][20] , \Term[4][19] , \Term[4][18] , 
        \Term[4][17] , \Term[4][16] , \Term[4][15] , \Term[4][14] , 
        \Term[4][13] , \Term[4][12] , \Term[4][11] , \Term[4][10] , 
        \Term[4][9] , \Term[4][8] , \Term[4][7] , \Term[4][6] , \Term[4][5] , 
        \Term[4][4] , \Term[4][3] , \Term[4][2] , \Term[4][1] , \Term[4][0] }), 
        .B({\Res[3][31] , \Res[3][30] , \Res[3][29] , \Res[3][28] , 
        \Res[3][27] , \Res[3][26] , \Res[3][25] , \Res[3][24] , \Res[3][23] , 
        \Res[3][22] , \Res[3][21] , \Res[3][20] , \Res[3][19] , \Res[3][18] , 
        \Res[3][17] , \Res[3][16] , \Res[3][15] , \Res[3][14] , \Res[3][13] , 
        \Res[3][12] , \Res[3][11] , \Res[3][10] , \Res[3][9] , \Res[3][8] , 
        \Res[3][7] , \Res[3][6] , \Res[3][5] , \Res[3][4] , \Res[3][3] , 
        \Res[3][2] , \Res[3][1] , \Res[3][0] }), .Ci(OP[4]), .S({\Res[4][31] , 
        \Res[4][30] , \Res[4][29] , \Res[4][28] , \Res[4][27] , \Res[4][26] , 
        \Res[4][25] , \Res[4][24] , \Res[4][23] , \Res[4][22] , \Res[4][21] , 
        \Res[4][20] , \Res[4][19] , \Res[4][18] , \Res[4][17] , \Res[4][16] , 
        \Res[4][15] , \Res[4][14] , \Res[4][13] , \Res[4][12] , \Res[4][11] , 
        \Res[4][10] , \Res[4][9] , \Res[4][8] , \Res[4][7] , \Res[4][6] , 
        \Res[4][5] , \Res[4][4] , \Res[4][3] , \Res[4][2] , \Res[4][1] , 
        \Res[4][0] }) );
  p4addgen_NB32_CW4_2 add_map_5 ( .A({\Term[5][31] , \Term[5][30] , 
        \Term[5][29] , \Term[5][28] , \Term[5][27] , \Term[5][26] , 
        \Term[5][25] , \Term[5][24] , \Term[5][23] , \Term[5][22] , 
        \Term[5][21] , \Term[5][20] , \Term[5][19] , \Term[5][18] , 
        \Term[5][17] , \Term[5][16] , \Term[5][15] , \Term[5][14] , 
        \Term[5][13] , \Term[5][12] , \Term[5][11] , \Term[5][10] , 
        \Term[5][9] , \Term[5][8] , \Term[5][7] , \Term[5][6] , \Term[5][5] , 
        \Term[5][4] , \Term[5][3] , \Term[5][2] , \Term[5][1] , \Term[5][0] }), 
        .B({\Res[4][31] , \Res[4][30] , \Res[4][29] , \Res[4][28] , 
        \Res[4][27] , \Res[4][26] , \Res[4][25] , \Res[4][24] , \Res[4][23] , 
        \Res[4][22] , \Res[4][21] , \Res[4][20] , \Res[4][19] , \Res[4][18] , 
        \Res[4][17] , \Res[4][16] , \Res[4][15] , \Res[4][14] , \Res[4][13] , 
        \Res[4][12] , \Res[4][11] , \Res[4][10] , \Res[4][9] , \Res[4][8] , 
        \Res[4][7] , \Res[4][6] , \Res[4][5] , \Res[4][4] , \Res[4][3] , 
        \Res[4][2] , \Res[4][1] , \Res[4][0] }), .Ci(OP[5]), .S({\Res[5][31] , 
        \Res[5][30] , \Res[5][29] , \Res[5][28] , \Res[5][27] , \Res[5][26] , 
        \Res[5][25] , \Res[5][24] , \Res[5][23] , \Res[5][22] , \Res[5][21] , 
        \Res[5][20] , \Res[5][19] , \Res[5][18] , \Res[5][17] , \Res[5][16] , 
        \Res[5][15] , \Res[5][14] , \Res[5][13] , \Res[5][12] , \Res[5][11] , 
        \Res[5][10] , \Res[5][9] , \Res[5][8] , \Res[5][7] , \Res[5][6] , 
        \Res[5][5] , \Res[5][4] , \Res[5][3] , \Res[5][2] , \Res[5][1] , 
        \Res[5][0] }) );
  p4addgen_NB32_CW4_1 add_map_6 ( .A({\Term[6][31] , \Term[6][30] , 
        \Term[6][29] , \Term[6][28] , \Term[6][27] , \Term[6][26] , 
        \Term[6][25] , \Term[6][24] , \Term[6][23] , \Term[6][22] , 
        \Term[6][21] , \Term[6][20] , \Term[6][19] , \Term[6][18] , 
        \Term[6][17] , \Term[6][16] , \Term[6][15] , \Term[6][14] , 
        \Term[6][13] , \Term[6][12] , \Term[6][11] , \Term[6][10] , 
        \Term[6][9] , \Term[6][8] , \Term[6][7] , \Term[6][6] , \Term[6][5] , 
        \Term[6][4] , \Term[6][3] , \Term[6][2] , \Term[6][1] , \Term[6][0] }), 
        .B({\Res[5][31] , \Res[5][30] , \Res[5][29] , \Res[5][28] , 
        \Res[5][27] , \Res[5][26] , \Res[5][25] , \Res[5][24] , \Res[5][23] , 
        \Res[5][22] , \Res[5][21] , \Res[5][20] , \Res[5][19] , \Res[5][18] , 
        \Res[5][17] , \Res[5][16] , \Res[5][15] , \Res[5][14] , \Res[5][13] , 
        \Res[5][12] , \Res[5][11] , \Res[5][10] , \Res[5][9] , \Res[5][8] , 
        \Res[5][7] , \Res[5][6] , \Res[5][5] , \Res[5][4] , \Res[5][3] , 
        \Res[5][2] , \Res[5][1] , \Res[5][0] }), .Ci(OP[6]), .S({\Res[6][31] , 
        \Res[6][30] , \Res[6][29] , \Res[6][28] , \Res[6][27] , \Res[6][26] , 
        \Res[6][25] , \Res[6][24] , \Res[6][23] , \Res[6][22] , \Res[6][21] , 
        \Res[6][20] , \Res[6][19] , \Res[6][18] , \Res[6][17] , \Res[6][16] , 
        \Res[6][15] , \Res[6][14] , \Res[6][13] , \Res[6][12] , \Res[6][11] , 
        \Res[6][10] , \Res[6][9] , \Res[6][8] , \Res[6][7] , \Res[6][6] , 
        \Res[6][5] , \Res[6][4] , \Res[6][3] , \Res[6][2] , \Res[6][1] , 
        \Res[6][0] }) );
  p4addgen_NB32_CW4_0 add_map_7 ( .A({\Term[7][31] , \Term[7][30] , 
        \Term[7][29] , \Term[7][28] , \Term[7][27] , \Term[7][26] , 
        \Term[7][25] , \Term[7][24] , \Term[7][23] , \Term[7][22] , 
        \Term[7][21] , \Term[7][20] , \Term[7][19] , \Term[7][18] , 
        \Term[7][17] , \Term[7][16] , \Term[7][15] , \Term[7][14] , 
        \Term[7][13] , \Term[7][12] , \Term[7][11] , \Term[7][10] , 
        \Term[7][9] , \Term[7][8] , \Term[7][7] , \Term[7][6] , \Term[7][5] , 
        \Term[7][4] , \Term[7][3] , \Term[7][2] , \Term[7][1] , \Term[7][0] }), 
        .B({\Res[6][31] , \Res[6][30] , \Res[6][29] , \Res[6][28] , 
        \Res[6][27] , \Res[6][26] , \Res[6][25] , \Res[6][24] , \Res[6][23] , 
        \Res[6][22] , \Res[6][21] , \Res[6][20] , \Res[6][19] , \Res[6][18] , 
        \Res[6][17] , \Res[6][16] , \Res[6][15] , \Res[6][14] , \Res[6][13] , 
        \Res[6][12] , \Res[6][11] , \Res[6][10] , \Res[6][9] , \Res[6][8] , 
        \Res[6][7] , \Res[6][6] , \Res[6][5] , \Res[6][4] , \Res[6][3] , 
        \Res[6][2] , \Res[6][1] , \Res[6][0] }), .Ci(OP[7]), .S(C) );
endmodule


module p4addgen_NB32_CW4_8 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [7:1] carry_sh;

  CLKBUF_X1 U1 ( .A(B[4]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(B[5]), .Z(n2) );
  BUF_X1 U3 ( .A(B[10]), .Z(n9) );
  CLKBUF_X1 U4 ( .A(B[3]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(B[7]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(B[13]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[9]), .Z(n6) );
  CLKBUF_X1 U8 ( .A(B[0]), .Z(n7) );
  CLKBUF_X1 U9 ( .A(B[12]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(A[0]), .Z(n10) );
  CLKBUF_X1 U11 ( .A(B[1]), .Z(n11) );
  CSTgen_CW4_NB32_8 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_8 carry_sel ( .A({A[31:1], n10}), .B({B[31:14], n5, n8, 
        B[11], n9, n6, B[8], n4, B[6], n2, n1, n3, B[2], n11, n7}), .Ci({
        carry_sh, Ci}), .S(S) );
endmodule


module MUX31_generic_NB32_0 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n7, n9, n10, n11, n12, n13, n14, n15, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n114, n8, n6, n5, n20, n19,
         n18, n113, n17, n16, n115;

  OAI221_X1 U2 ( .B1(n14), .B2(n44), .C1(n1), .C2(n43), .A(n42), .ZN(Y[8]) );
  OAI221_X1 U3 ( .B1(n15), .B2(n107), .C1(n12), .C2(n106), .A(n105), .ZN(Y[29]) );
  OAI221_X1 U11 ( .B1(n41), .B2(n14), .C1(n1), .C2(n40), .A(n39), .ZN(Y[7]) );
  CLKBUF_X1 U12 ( .A(n11), .Z(n1) );
  OAI221_X1 U13 ( .B1(n14), .B2(n26), .C1(n10), .C2(n25), .A(n24), .ZN(Y[2])
         );
  CLKBUF_X1 U14 ( .A(n14), .Z(n2) );
  OAI221_X1 U15 ( .B1(n15), .B2(n62), .C1(n12), .C2(n61), .A(n60), .ZN(Y[14])
         );
  OAI221_X1 U16 ( .B1(n50), .B2(n15), .C1(n10), .C2(n49), .A(n48), .ZN(Y[10])
         );
  OAI221_X1 U17 ( .B1(n14), .B2(n95), .C1(n12), .C2(n94), .A(n93), .ZN(Y[25])
         );
  OAI221_X1 U18 ( .B1(n86), .B2(n14), .C1(n10), .C2(n85), .A(n84), .ZN(Y[22])
         );
  OAI221_X1 U19 ( .B1(n14), .B2(n89), .C1(n12), .C2(n88), .A(n87), .ZN(Y[23])
         );
  OAI221_X1 U20 ( .B1(n15), .B2(n98), .C1(n12), .C2(n97), .A(n96), .ZN(Y[26])
         );
  OAI221_X1 U21 ( .B1(n14), .B2(n65), .C1(n12), .C2(n64), .A(n63), .ZN(Y[15])
         );
  OAI221_X1 U23 ( .B1(n14), .B2(n104), .C1(n10), .C2(n103), .A(n102), .ZN(
        Y[28]) );
  OAI221_X1 U24 ( .B1(n15), .B2(n74), .C1(n12), .C2(n73), .A(n72), .ZN(Y[18])
         );
  OAI221_X1 U25 ( .B1(n15), .B2(n83), .C1(n10), .C2(n82), .A(n81), .ZN(Y[21])
         );
  OAI221_X1 U27 ( .B1(n15), .B2(n38), .C1(n10), .C2(n37), .A(n36), .ZN(Y[6])
         );
  OAI221_X1 U28 ( .B1(n14), .B2(n71), .C1(n10), .C2(n70), .A(n69), .ZN(Y[17])
         );
  OAI221_X1 U29 ( .B1(n14), .B2(n35), .C1(n10), .C2(n34), .A(n33), .ZN(Y[5])
         );
  OAI221_X4 U32 ( .B1(n15), .B2(n32), .C1(n12), .C2(n31), .A(n30), .ZN(Y[4])
         );
  OAI221_X1 U33 ( .B1(n29), .B2(n13), .C1(n10), .C2(n28), .A(n27), .ZN(Y[3])
         );
  OAI221_X1 U35 ( .B1(n15), .B2(n114), .C1(n1), .C2(n112), .A(n111), .ZN(Y[31]) );
  OAI221_X1 U36 ( .B1(n14), .B2(n101), .C1(n10), .C2(n100), .A(n99), .ZN(Y[27]) );
  OAI221_X1 U37 ( .B1(n2), .B2(n110), .C1(n12), .C2(n109), .A(n108), .ZN(Y[30]) );
  OAI221_X1 U38 ( .B1(n14), .B2(n56), .C1(n10), .C2(n55), .A(n54), .ZN(Y[12])
         );
  OAI221_X4 U40 ( .B1(n47), .B2(n13), .C1(n11), .C2(n46), .A(n45), .ZN(Y[9])
         );
  OAI221_X4 U42 ( .B1(n13), .B2(n23), .C1(n11), .C2(n22), .A(n21), .ZN(Y[1])
         );
  INV_X1 U52 ( .A(C[1]), .ZN(n23) );
  INV_X1 U53 ( .A(A[1]), .ZN(n22) );
  INV_X1 U55 ( .A(C[2]), .ZN(n26) );
  INV_X1 U56 ( .A(A[2]), .ZN(n25) );
  NAND2_X1 U57 ( .A1(B[2]), .A2(n7), .ZN(n24) );
  INV_X1 U58 ( .A(C[3]), .ZN(n29) );
  INV_X1 U59 ( .A(A[3]), .ZN(n28) );
  NAND2_X1 U60 ( .A1(n7), .A2(B[3]), .ZN(n27) );
  INV_X1 U61 ( .A(C[4]), .ZN(n32) );
  INV_X1 U62 ( .A(A[4]), .ZN(n31) );
  NAND2_X1 U63 ( .A1(B[4]), .A2(n3), .ZN(n30) );
  INV_X1 U64 ( .A(C[5]), .ZN(n35) );
  INV_X1 U65 ( .A(A[5]), .ZN(n34) );
  NAND2_X1 U66 ( .A1(n4), .A2(B[5]), .ZN(n33) );
  INV_X1 U67 ( .A(C[6]), .ZN(n38) );
  INV_X1 U68 ( .A(A[6]), .ZN(n37) );
  NAND2_X1 U69 ( .A1(B[6]), .A2(n3), .ZN(n36) );
  INV_X1 U70 ( .A(C[7]), .ZN(n41) );
  INV_X1 U71 ( .A(A[7]), .ZN(n40) );
  NAND2_X1 U72 ( .A1(B[7]), .A2(n3), .ZN(n39) );
  INV_X1 U73 ( .A(C[8]), .ZN(n44) );
  INV_X1 U74 ( .A(A[8]), .ZN(n43) );
  NAND2_X1 U75 ( .A1(B[8]), .A2(n3), .ZN(n42) );
  INV_X1 U76 ( .A(C[9]), .ZN(n47) );
  INV_X1 U77 ( .A(A[9]), .ZN(n46) );
  INV_X1 U79 ( .A(C[10]), .ZN(n50) );
  INV_X1 U80 ( .A(A[10]), .ZN(n49) );
  NAND2_X1 U81 ( .A1(B[10]), .A2(n3), .ZN(n48) );
  INV_X1 U82 ( .A(C[11]), .ZN(n53) );
  INV_X1 U83 ( .A(A[11]), .ZN(n52) );
  NAND2_X1 U84 ( .A1(B[11]), .A2(n7), .ZN(n51) );
  INV_X1 U85 ( .A(C[12]), .ZN(n56) );
  INV_X1 U86 ( .A(A[12]), .ZN(n55) );
  NAND2_X1 U87 ( .A1(B[12]), .A2(n9), .ZN(n54) );
  INV_X1 U88 ( .A(C[13]), .ZN(n59) );
  INV_X1 U89 ( .A(A[13]), .ZN(n58) );
  NAND2_X1 U90 ( .A1(B[13]), .A2(n4), .ZN(n57) );
  INV_X1 U91 ( .A(C[14]), .ZN(n62) );
  INV_X1 U92 ( .A(A[14]), .ZN(n61) );
  NAND2_X1 U93 ( .A1(B[14]), .A2(n7), .ZN(n60) );
  INV_X1 U94 ( .A(C[15]), .ZN(n65) );
  INV_X1 U95 ( .A(A[15]), .ZN(n64) );
  NAND2_X1 U96 ( .A1(B[15]), .A2(n7), .ZN(n63) );
  INV_X1 U97 ( .A(C[16]), .ZN(n68) );
  INV_X1 U98 ( .A(A[16]), .ZN(n67) );
  NAND2_X1 U99 ( .A1(B[16]), .A2(n4), .ZN(n66) );
  OAI221_X1 U100 ( .B1(n14), .B2(n68), .C1(n10), .C2(n67), .A(n66), .ZN(Y[16])
         );
  INV_X1 U101 ( .A(C[17]), .ZN(n71) );
  INV_X1 U102 ( .A(A[17]), .ZN(n70) );
  NAND2_X1 U103 ( .A1(B[17]), .A2(n7), .ZN(n69) );
  INV_X1 U104 ( .A(C[18]), .ZN(n74) );
  INV_X1 U105 ( .A(A[18]), .ZN(n73) );
  NAND2_X1 U106 ( .A1(B[18]), .A2(n9), .ZN(n72) );
  INV_X1 U107 ( .A(C[19]), .ZN(n77) );
  INV_X1 U108 ( .A(A[19]), .ZN(n76) );
  NAND2_X1 U109 ( .A1(B[19]), .A2(n3), .ZN(n75) );
  OAI221_X1 U110 ( .B1(n15), .B2(n77), .C1(n12), .C2(n76), .A(n75), .ZN(Y[19])
         );
  INV_X1 U111 ( .A(C[20]), .ZN(n80) );
  INV_X1 U112 ( .A(A[20]), .ZN(n79) );
  NAND2_X1 U113 ( .A1(B[20]), .A2(n7), .ZN(n78) );
  OAI221_X1 U114 ( .B1(n15), .B2(n80), .C1(n12), .C2(n79), .A(n78), .ZN(Y[20])
         );
  INV_X1 U115 ( .A(C[21]), .ZN(n83) );
  INV_X1 U116 ( .A(A[21]), .ZN(n82) );
  NAND2_X1 U117 ( .A1(n7), .A2(B[21]), .ZN(n81) );
  INV_X1 U118 ( .A(C[22]), .ZN(n86) );
  INV_X1 U119 ( .A(A[22]), .ZN(n85) );
  NAND2_X1 U120 ( .A1(B[22]), .A2(n9), .ZN(n84) );
  INV_X1 U121 ( .A(C[23]), .ZN(n89) );
  INV_X1 U122 ( .A(A[23]), .ZN(n88) );
  NAND2_X1 U123 ( .A1(B[23]), .A2(n7), .ZN(n87) );
  INV_X1 U124 ( .A(C[24]), .ZN(n92) );
  INV_X1 U125 ( .A(A[24]), .ZN(n91) );
  NAND2_X1 U126 ( .A1(B[24]), .A2(n3), .ZN(n90) );
  OAI221_X1 U127 ( .B1(n15), .B2(n92), .C1(n12), .C2(n91), .A(n90), .ZN(Y[24])
         );
  INV_X1 U128 ( .A(C[25]), .ZN(n95) );
  INV_X1 U129 ( .A(A[25]), .ZN(n94) );
  NAND2_X1 U130 ( .A1(B[25]), .A2(n4), .ZN(n93) );
  INV_X1 U131 ( .A(C[26]), .ZN(n98) );
  INV_X1 U132 ( .A(A[26]), .ZN(n97) );
  NAND2_X1 U133 ( .A1(B[26]), .A2(n7), .ZN(n96) );
  INV_X1 U134 ( .A(C[27]), .ZN(n101) );
  INV_X1 U135 ( .A(A[27]), .ZN(n100) );
  NAND2_X1 U136 ( .A1(B[27]), .A2(n3), .ZN(n99) );
  INV_X1 U137 ( .A(C[28]), .ZN(n104) );
  INV_X1 U138 ( .A(A[28]), .ZN(n103) );
  NAND2_X1 U139 ( .A1(B[28]), .A2(n4), .ZN(n102) );
  INV_X1 U140 ( .A(C[29]), .ZN(n107) );
  INV_X1 U141 ( .A(A[29]), .ZN(n106) );
  NAND2_X1 U142 ( .A1(B[29]), .A2(n7), .ZN(n105) );
  INV_X1 U143 ( .A(C[30]), .ZN(n110) );
  INV_X1 U144 ( .A(A[30]), .ZN(n109) );
  NAND2_X1 U145 ( .A1(n3), .A2(B[30]), .ZN(n108) );
  INV_X1 U146 ( .A(C[31]), .ZN(n114) );
  INV_X1 U147 ( .A(A[31]), .ZN(n112) );
  NAND2_X1 U148 ( .A1(B[31]), .A2(n4), .ZN(n111) );
  CLKBUF_X3 U45 ( .A(n113), .Z(n10) );
  CLKBUF_X3 U34 ( .A(n113), .Z(n12) );
  AND2_X2 U39 ( .A1(n5), .A2(n6), .ZN(n7) );
  AND2_X1 U8 ( .A1(n5), .A2(n6), .ZN(n3) );
  NAND2_X1 U54 ( .A1(B[1]), .A2(n8), .ZN(n21) );
  NAND2_X1 U78 ( .A1(n4), .A2(B[9]), .ZN(n45) );
  INV_X1 U47 ( .A(C[0]), .ZN(n20) );
  INV_X1 U49 ( .A(A[0]), .ZN(n19) );
  NAND2_X1 U50 ( .A1(B[0]), .A2(n8), .ZN(n18) );
  OAI221_X1 U51 ( .B1(n13), .B2(n20), .C1(n11), .C2(n19), .A(n18), .ZN(Y[0])
         );
  BUF_X1 U7 ( .A(SEL[0]), .Z(n5) );
  INV_X1 U48 ( .A(SEL[1]), .ZN(n17) );
  INV_X1 U41 ( .A(SEL[1]), .ZN(n6) );
  NAND2_X1 U44 ( .A1(n17), .A2(n16), .ZN(n113) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n16) );
  BUF_X2 U22 ( .A(n115), .Z(n13) );
  CLKBUF_X3 U10 ( .A(n115), .Z(n15) );
  CLKBUF_X3 U9 ( .A(n115), .Z(n14) );
  NAND2_X1 U43 ( .A1(SEL[1]), .A2(n16), .ZN(n115) );
  OAI221_X1 U4 ( .B1(n15), .B2(n59), .C1(n12), .C2(n58), .A(n57), .ZN(Y[13])
         );
  OAI221_X1 U5 ( .B1(n53), .B2(n13), .C1(n11), .C2(n52), .A(n51), .ZN(Y[11])
         );
  BUF_X2 U6 ( .A(n113), .Z(n11) );
  AND2_X2 U26 ( .A1(n5), .A2(n6), .ZN(n4) );
  AND2_X1 U30 ( .A1(n5), .A2(n17), .ZN(n8) );
  BUF_X1 U31 ( .A(n4), .Z(n9) );
endmodule


module MUX31_generic_NB32_1 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n146;

  OAI221_X4 U2 ( .B1(n15), .B2(n33), .C1(n12), .C2(n32), .A(n31), .ZN(Y[4]) );
  OAI221_X4 U3 ( .B1(n14), .B2(n63), .C1(n11), .C2(n62), .A(n61), .ZN(Y[14])
         );
  NAND3_X2 U4 ( .A1(n2), .A2(n3), .A3(n64), .ZN(Y[15]) );
  AND2_X1 U5 ( .A1(SEL[0]), .A2(n1), .ZN(n7) );
  OAI221_X4 U6 ( .B1(n13), .B2(n102), .C1(n10), .C2(n101), .A(n100), .ZN(Y[27]) );
  CLKBUF_X3 U7 ( .A(n114), .Z(n10) );
  CLKBUF_X3 U8 ( .A(n116), .Z(n13) );
  INV_X1 U9 ( .A(SEL[1]), .ZN(n1) );
  OAI221_X4 U10 ( .B1(n15), .B2(n42), .C1(n12), .C2(n41), .A(n40), .ZN(Y[7])
         );
  OR2_X1 U11 ( .A1(n14), .A2(n66), .ZN(n2) );
  OR2_X1 U12 ( .A1(n11), .A2(n65), .ZN(n3) );
  BUF_X2 U13 ( .A(n116), .Z(n14) );
  OR2_X1 U14 ( .A1(n14), .A2(n54), .ZN(n4) );
  OR2_X1 U15 ( .A1(n11), .A2(n53), .ZN(n5) );
  NAND3_X1 U16 ( .A1(n4), .A2(n5), .A3(n52), .ZN(Y[11]) );
  OAI221_X4 U17 ( .B1(n15), .B2(n30), .C1(n12), .C2(n29), .A(n28), .ZN(Y[3])
         );
  OAI221_X4 U18 ( .B1(n13), .B2(n90), .C1(n10), .C2(n89), .A(n88), .ZN(Y[23])
         );
  OAI221_X4 U19 ( .B1(n13), .B2(n81), .C1(n10), .C2(n80), .A(n79), .ZN(Y[20])
         );
  OAI221_X4 U20 ( .B1(n13), .B2(n93), .C1(n10), .C2(n92), .A(n91), .ZN(Y[24])
         );
  OAI221_X4 U21 ( .B1(n14), .B2(n78), .C1(n11), .C2(n77), .A(n76), .ZN(Y[19])
         );
  OAI221_X4 U22 ( .B1(n13), .B2(n108), .C1(n10), .C2(n107), .A(n106), .ZN(
        Y[29]) );
  OAI221_X4 U23 ( .B1(n13), .B2(n87), .C1(n10), .C2(n86), .A(n85), .ZN(Y[22])
         );
  OAI221_X4 U24 ( .B1(n14), .B2(n69), .C1(n11), .C2(n68), .A(n67), .ZN(Y[16])
         );
  OAI221_X4 U25 ( .B1(n13), .B2(n99), .C1(n10), .C2(n98), .A(n97), .ZN(Y[26])
         );
  OAI221_X4 U26 ( .B1(n14), .B2(n75), .C1(n11), .C2(n74), .A(n73), .ZN(Y[18])
         );
  OAI221_X4 U27 ( .B1(n13), .B2(n84), .C1(n10), .C2(n83), .A(n82), .ZN(Y[21])
         );
  OAI221_X4 U28 ( .B1(n13), .B2(n105), .C1(n10), .C2(n104), .A(n103), .ZN(
        Y[28]) );
  OAI221_X4 U29 ( .B1(n14), .B2(n72), .C1(n11), .C2(n71), .A(n70), .ZN(Y[17])
         );
  OAI221_X4 U30 ( .B1(n13), .B2(n96), .C1(n10), .C2(n95), .A(n94), .ZN(Y[25])
         );
  AND2_X2 U31 ( .A1(SEL[0]), .A2(n18), .ZN(n6) );
  BUF_X2 U32 ( .A(n114), .Z(n11) );
  BUF_X2 U33 ( .A(n114), .Z(n12) );
  BUF_X2 U34 ( .A(n116), .Z(n15) );
  NAND2_X1 U35 ( .A1(n17), .A2(SEL[1]), .ZN(n116) );
  BUF_X2 U37 ( .A(n7), .Z(n9) );
  BUF_X1 U38 ( .A(n146), .Z(Y[2]) );
  NAND2_X1 U39 ( .A1(n17), .A2(n18), .ZN(n114) );
  INV_X1 U40 ( .A(SEL[0]), .ZN(n17) );
  INV_X1 U41 ( .A(C[0]), .ZN(n21) );
  INV_X1 U42 ( .A(SEL[1]), .ZN(n18) );
  INV_X1 U43 ( .A(A[0]), .ZN(n20) );
  NAND2_X1 U44 ( .A1(n9), .A2(B[0]), .ZN(n19) );
  OAI221_X1 U45 ( .B1(n15), .B2(n21), .C1(n12), .C2(n20), .A(n19), .ZN(Y[0])
         );
  INV_X1 U46 ( .A(C[1]), .ZN(n24) );
  INV_X1 U47 ( .A(A[1]), .ZN(n23) );
  NAND2_X1 U48 ( .A1(B[1]), .A2(n9), .ZN(n22) );
  OAI221_X1 U49 ( .B1(n15), .B2(n24), .C1(n12), .C2(n23), .A(n22), .ZN(Y[1])
         );
  INV_X1 U50 ( .A(C[2]), .ZN(n27) );
  INV_X1 U51 ( .A(A[2]), .ZN(n26) );
  NAND2_X1 U52 ( .A1(B[2]), .A2(n9), .ZN(n25) );
  OAI221_X1 U53 ( .B1(n15), .B2(n27), .C1(n12), .C2(n26), .A(n25), .ZN(n146)
         );
  INV_X1 U54 ( .A(C[3]), .ZN(n30) );
  INV_X1 U55 ( .A(A[3]), .ZN(n29) );
  NAND2_X1 U56 ( .A1(B[3]), .A2(n8), .ZN(n28) );
  INV_X1 U57 ( .A(C[4]), .ZN(n33) );
  INV_X1 U58 ( .A(A[4]), .ZN(n32) );
  NAND2_X1 U59 ( .A1(B[4]), .A2(n6), .ZN(n31) );
  INV_X1 U60 ( .A(C[5]), .ZN(n36) );
  INV_X1 U61 ( .A(A[5]), .ZN(n35) );
  NAND2_X1 U62 ( .A1(B[5]), .A2(n8), .ZN(n34) );
  OAI221_X1 U63 ( .B1(n15), .B2(n36), .C1(n12), .C2(n35), .A(n34), .ZN(Y[5])
         );
  INV_X1 U64 ( .A(C[6]), .ZN(n39) );
  INV_X1 U65 ( .A(A[6]), .ZN(n38) );
  NAND2_X1 U66 ( .A1(B[6]), .A2(n9), .ZN(n37) );
  OAI221_X1 U67 ( .B1(n15), .B2(n39), .C1(n12), .C2(n38), .A(n37), .ZN(Y[6])
         );
  INV_X1 U68 ( .A(C[7]), .ZN(n42) );
  INV_X1 U69 ( .A(A[7]), .ZN(n41) );
  NAND2_X1 U70 ( .A1(B[7]), .A2(n8), .ZN(n40) );
  INV_X1 U71 ( .A(C[8]), .ZN(n45) );
  INV_X1 U72 ( .A(A[8]), .ZN(n44) );
  NAND2_X1 U73 ( .A1(B[8]), .A2(n8), .ZN(n43) );
  OAI221_X1 U74 ( .B1(n14), .B2(n45), .C1(n11), .C2(n44), .A(n43), .ZN(Y[8])
         );
  INV_X1 U75 ( .A(C[9]), .ZN(n48) );
  INV_X1 U76 ( .A(A[9]), .ZN(n47) );
  NAND2_X1 U77 ( .A1(B[9]), .A2(n9), .ZN(n46) );
  OAI221_X1 U78 ( .B1(n14), .B2(n48), .C1(n11), .C2(n47), .A(n46), .ZN(Y[9])
         );
  INV_X1 U79 ( .A(C[10]), .ZN(n51) );
  INV_X1 U80 ( .A(A[10]), .ZN(n50) );
  NAND2_X1 U81 ( .A1(B[10]), .A2(n8), .ZN(n49) );
  OAI221_X1 U82 ( .B1(n14), .B2(n51), .C1(n11), .C2(n50), .A(n49), .ZN(Y[10])
         );
  INV_X1 U83 ( .A(C[11]), .ZN(n54) );
  INV_X1 U84 ( .A(A[11]), .ZN(n53) );
  NAND2_X1 U85 ( .A1(B[11]), .A2(n8), .ZN(n52) );
  INV_X1 U86 ( .A(C[12]), .ZN(n57) );
  INV_X1 U87 ( .A(A[12]), .ZN(n56) );
  NAND2_X1 U88 ( .A1(B[12]), .A2(n6), .ZN(n55) );
  OAI221_X1 U89 ( .B1(n14), .B2(n57), .C1(n11), .C2(n56), .A(n55), .ZN(Y[12])
         );
  INV_X1 U90 ( .A(C[13]), .ZN(n60) );
  INV_X1 U91 ( .A(A[13]), .ZN(n59) );
  NAND2_X1 U92 ( .A1(B[13]), .A2(n9), .ZN(n58) );
  OAI221_X1 U93 ( .B1(n14), .B2(n60), .C1(n11), .C2(n59), .A(n58), .ZN(Y[13])
         );
  INV_X1 U94 ( .A(C[14]), .ZN(n63) );
  INV_X1 U95 ( .A(A[14]), .ZN(n62) );
  NAND2_X1 U96 ( .A1(B[14]), .A2(n6), .ZN(n61) );
  INV_X1 U97 ( .A(C[15]), .ZN(n66) );
  INV_X1 U98 ( .A(A[15]), .ZN(n65) );
  NAND2_X1 U99 ( .A1(B[15]), .A2(n8), .ZN(n64) );
  INV_X1 U100 ( .A(C[16]), .ZN(n69) );
  INV_X1 U101 ( .A(A[16]), .ZN(n68) );
  NAND2_X1 U102 ( .A1(B[16]), .A2(n8), .ZN(n67) );
  INV_X1 U103 ( .A(C[17]), .ZN(n72) );
  INV_X1 U104 ( .A(A[17]), .ZN(n71) );
  NAND2_X1 U105 ( .A1(B[17]), .A2(n6), .ZN(n70) );
  INV_X1 U106 ( .A(C[18]), .ZN(n75) );
  INV_X1 U107 ( .A(A[18]), .ZN(n74) );
  NAND2_X1 U108 ( .A1(B[18]), .A2(n8), .ZN(n73) );
  INV_X1 U109 ( .A(C[19]), .ZN(n78) );
  INV_X1 U110 ( .A(A[19]), .ZN(n77) );
  NAND2_X1 U111 ( .A1(B[19]), .A2(n6), .ZN(n76) );
  INV_X1 U112 ( .A(C[20]), .ZN(n81) );
  INV_X1 U113 ( .A(A[20]), .ZN(n80) );
  NAND2_X1 U114 ( .A1(B[20]), .A2(n6), .ZN(n79) );
  INV_X1 U115 ( .A(C[21]), .ZN(n84) );
  INV_X1 U116 ( .A(A[21]), .ZN(n83) );
  NAND2_X1 U117 ( .A1(B[21]), .A2(n6), .ZN(n82) );
  INV_X1 U118 ( .A(C[22]), .ZN(n87) );
  INV_X1 U119 ( .A(A[22]), .ZN(n86) );
  NAND2_X1 U120 ( .A1(B[22]), .A2(n6), .ZN(n85) );
  INV_X1 U121 ( .A(C[23]), .ZN(n90) );
  INV_X1 U122 ( .A(A[23]), .ZN(n89) );
  NAND2_X1 U123 ( .A1(B[23]), .A2(n6), .ZN(n88) );
  INV_X1 U124 ( .A(C[24]), .ZN(n93) );
  INV_X1 U125 ( .A(A[24]), .ZN(n92) );
  NAND2_X1 U126 ( .A1(B[24]), .A2(n6), .ZN(n91) );
  INV_X1 U127 ( .A(C[25]), .ZN(n96) );
  INV_X1 U128 ( .A(A[25]), .ZN(n95) );
  NAND2_X1 U129 ( .A1(B[25]), .A2(n8), .ZN(n94) );
  INV_X1 U130 ( .A(C[26]), .ZN(n99) );
  INV_X1 U131 ( .A(A[26]), .ZN(n98) );
  NAND2_X1 U132 ( .A1(B[26]), .A2(n6), .ZN(n97) );
  INV_X1 U133 ( .A(C[27]), .ZN(n102) );
  INV_X1 U134 ( .A(A[27]), .ZN(n101) );
  NAND2_X1 U135 ( .A1(B[27]), .A2(n6), .ZN(n100) );
  INV_X1 U136 ( .A(C[28]), .ZN(n105) );
  INV_X1 U137 ( .A(A[28]), .ZN(n104) );
  NAND2_X1 U138 ( .A1(B[28]), .A2(n8), .ZN(n103) );
  INV_X1 U139 ( .A(C[29]), .ZN(n108) );
  INV_X1 U140 ( .A(A[29]), .ZN(n107) );
  NAND2_X1 U141 ( .A1(B[29]), .A2(n8), .ZN(n106) );
  INV_X1 U142 ( .A(C[30]), .ZN(n111) );
  INV_X1 U143 ( .A(A[30]), .ZN(n110) );
  NAND2_X1 U144 ( .A1(B[30]), .A2(n6), .ZN(n109) );
  OAI221_X1 U145 ( .B1(n13), .B2(n111), .C1(n10), .C2(n110), .A(n109), .ZN(
        Y[30]) );
  INV_X1 U146 ( .A(C[31]), .ZN(n115) );
  INV_X1 U147 ( .A(A[31]), .ZN(n113) );
  NAND2_X1 U148 ( .A1(B[31]), .A2(n6), .ZN(n112) );
  OAI221_X1 U149 ( .B1(n13), .B2(n115), .C1(n10), .C2(n113), .A(n112), .ZN(
        Y[31]) );
  CLKBUF_X3 U36 ( .A(n7), .Z(n8) );
endmodule


module MUX21_generic_NB32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  CLKBUF_X1 U1 ( .A(SEL), .Z(n3) );
  CLKBUF_X3 U2 ( .A(SEL), .Z(n1) );
  CLKBUF_X3 U3 ( .A(SEL), .Z(n2) );
  MUX2_X1 U4 ( .A(B[0]), .B(A[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(B[1]), .B(A[1]), .S(n1), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(B[2]), .B(A[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U7 ( .A(B[3]), .B(A[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U8 ( .A(B[4]), .B(A[4]), .S(n1), .Z(Y[4]) );
  MUX2_X1 U9 ( .A(B[5]), .B(A[5]), .S(n1), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(B[6]), .B(A[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(B[7]), .B(A[7]), .S(n1), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(B[8]), .B(A[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(B[9]), .B(A[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(B[10]), .B(A[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(B[11]), .B(A[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(B[12]), .B(A[12]), .S(n2), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(B[13]), .B(A[13]), .S(n2), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(B[14]), .B(A[14]), .S(n2), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(B[15]), .B(A[15]), .S(n2), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(B[16]), .B(A[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(B[17]), .B(A[17]), .S(n2), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(B[18]), .B(A[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(B[19]), .B(A[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(B[20]), .B(A[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(B[21]), .B(A[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(B[22]), .B(A[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(B[23]), .B(A[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(B[24]), .B(A[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(B[25]), .B(A[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(B[26]), .B(A[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(B[27]), .B(A[27]), .S(n3), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(B[28]), .B(A[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(B[29]), .B(A[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(B[30]), .B(A[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(B[31]), .B(A[31]), .S(n3), .Z(Y[31]) );
endmodule


module MUX21_generic_NB32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  CLKBUF_X1 U1 ( .A(SEL), .Z(n3) );
  BUF_X2 U2 ( .A(SEL), .Z(n2) );
  CLKBUF_X3 U3 ( .A(SEL), .Z(n1) );
  MUX2_X1 U4 ( .A(B[0]), .B(A[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(B[1]), .B(A[1]), .S(n1), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(B[2]), .B(A[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U7 ( .A(B[3]), .B(A[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U8 ( .A(B[4]), .B(A[4]), .S(n1), .Z(Y[4]) );
  MUX2_X1 U9 ( .A(B[5]), .B(A[5]), .S(n1), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(B[6]), .B(A[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(B[7]), .B(A[7]), .S(n1), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(B[8]), .B(A[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(B[9]), .B(A[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(B[10]), .B(A[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(B[11]), .B(A[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(B[12]), .B(A[12]), .S(n2), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(B[13]), .B(A[13]), .S(n2), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(B[14]), .B(A[14]), .S(n2), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(B[15]), .B(A[15]), .S(n2), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(B[16]), .B(A[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(B[17]), .B(A[17]), .S(n2), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(B[18]), .B(A[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(B[19]), .B(A[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(B[20]), .B(A[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(B[21]), .B(A[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(B[22]), .B(A[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(B[23]), .B(A[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(B[24]), .B(A[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(B[25]), .B(A[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(B[26]), .B(A[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(B[27]), .B(A[27]), .S(n3), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(B[28]), .B(A[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(B[29]), .B(A[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(B[30]), .B(A[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(B[31]), .B(A[31]), .S(n3), .Z(Y[31]) );
endmodule


module FD_INJ_NB5_0 ( CK, RESET, INJ_ZERO, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, INJ_ZERO;

  wire   [4:0] TMP_D;

  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  SDFFR_X1 \Q_reg[1]  ( .D(1'b0), .SI(INJ_ZERO), .SE(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  SDFFR_X1 \Q_reg[2]  ( .D(1'b0), .SI(INJ_ZERO), .SE(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  AND2_X1 U5 ( .A1(D[3]), .A2(INJ_ZERO), .ZN(TMP_D[3]) );
  AND2_X1 U6 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U7 ( .A1(INJ_ZERO), .A2(D[4]), .ZN(TMP_D[4]) );
endmodule


module FD_INJ_NB5_1 ( CK, RESET, INJ_ZERO, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, INJ_ZERO;

  wire   [4:0] TMP_D;

  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  SDFFR_X1 \Q_reg[2]  ( .D(1'b0), .SI(INJ_ZERO), .SE(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  AND2_X1 U4 ( .A1(INJ_ZERO), .A2(D[4]), .ZN(TMP_D[4]) );
  AND2_X1 U5 ( .A1(D[3]), .A2(INJ_ZERO), .ZN(TMP_D[3]) );
  AND2_X1 U6 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U7 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
endmodule


module FD_INJ_NB5_2 ( CK, RESET, INJ_ZERO, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, INJ_ZERO;

  wire   [4:0] TMP_D;

  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[4]), .ZN(TMP_D[4]) );
  AND2_X1 U4 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U5 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U6 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
  AND2_X1 U7 ( .A1(D[3]), .A2(INJ_ZERO), .ZN(TMP_D[3]) );
endmodule


module MUX21_generic_NB5_0 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;
  wire   n8, n9, n10, n11, n12, n13;

  INV_X1 U1 ( .A(n8), .ZN(Y[4]) );
  AOI22_X1 U2 ( .A1(SEL), .A2(A[4]), .B1(B[4]), .B2(n9), .ZN(n8) );
  INV_X1 U3 ( .A(n13), .ZN(Y[0]) );
  AOI22_X1 U4 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n9), .ZN(n13) );
  INV_X1 U5 ( .A(n12), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n9), .ZN(n12) );
  INV_X1 U7 ( .A(n11), .ZN(Y[2]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n9), .ZN(n11) );
  INV_X1 U9 ( .A(n10), .ZN(Y[3]) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(SEL), .B1(B[3]), .B2(n9), .ZN(n10) );
  INV_X1 U11 ( .A(SEL), .ZN(n9) );
endmodule


module FD_INJ_NB32_0 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n1, n34, n35, n36;
  wire   [31:0] TMP_D;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n36), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n36), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n36), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n36), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n36), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n36), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n36), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n36), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n35), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n35), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n35), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n35), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n35), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n35), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n35), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n35), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n35), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n35), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n35), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n35), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n34), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n34), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n34), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n34), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n34), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n34), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n34), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n34), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n34), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n34), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n34), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n34), .Q(Q[0]) );
  CLKBUF_X1 U3 ( .A(INJ_ZERO), .Z(n1) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
  BUF_X1 U6 ( .A(RESET), .Z(n36) );
  AND2_X1 U7 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U8 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U9 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
  AND2_X1 U10 ( .A1(D[10]), .A2(INJ_ZERO), .ZN(TMP_D[10]) );
  AND2_X1 U11 ( .A1(D[11]), .A2(INJ_ZERO), .ZN(TMP_D[11]) );
  AND2_X1 U12 ( .A1(D[12]), .A2(INJ_ZERO), .ZN(TMP_D[12]) );
  AND2_X1 U13 ( .A1(D[13]), .A2(INJ_ZERO), .ZN(TMP_D[13]) );
  AND2_X1 U14 ( .A1(D[14]), .A2(INJ_ZERO), .ZN(TMP_D[14]) );
  AND2_X1 U15 ( .A1(D[15]), .A2(n1), .ZN(TMP_D[15]) );
  AND2_X1 U16 ( .A1(D[16]), .A2(n1), .ZN(TMP_D[16]) );
  AND2_X1 U17 ( .A1(D[17]), .A2(n1), .ZN(TMP_D[17]) );
  AND2_X1 U18 ( .A1(D[18]), .A2(n1), .ZN(TMP_D[18]) );
  AND2_X1 U19 ( .A1(D[19]), .A2(INJ_ZERO), .ZN(TMP_D[19]) );
  AND2_X1 U20 ( .A1(D[20]), .A2(INJ_ZERO), .ZN(TMP_D[20]) );
  AND2_X1 U21 ( .A1(D[21]), .A2(INJ_ZERO), .ZN(TMP_D[21]) );
  AND2_X1 U22 ( .A1(D[22]), .A2(INJ_ZERO), .ZN(TMP_D[22]) );
  AND2_X1 U23 ( .A1(D[23]), .A2(INJ_ZERO), .ZN(TMP_D[23]) );
  AND2_X1 U24 ( .A1(D[24]), .A2(INJ_ZERO), .ZN(TMP_D[24]) );
  AND2_X1 U25 ( .A1(D[25]), .A2(INJ_ZERO), .ZN(TMP_D[25]) );
  AND2_X1 U26 ( .A1(D[26]), .A2(INJ_ZERO), .ZN(TMP_D[26]) );
  AND2_X1 U27 ( .A1(D[27]), .A2(INJ_ZERO), .ZN(TMP_D[27]) );
  AND2_X1 U28 ( .A1(D[28]), .A2(INJ_ZERO), .ZN(TMP_D[28]) );
  AND2_X1 U29 ( .A1(D[29]), .A2(INJ_ZERO), .ZN(TMP_D[29]) );
  AND2_X1 U30 ( .A1(D[30]), .A2(INJ_ZERO), .ZN(TMP_D[30]) );
  AND2_X1 U31 ( .A1(n1), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U32 ( .A1(D[3]), .A2(n1), .ZN(TMP_D[3]) );
  AND2_X1 U33 ( .A1(D[4]), .A2(n1), .ZN(TMP_D[4]) );
  AND2_X1 U34 ( .A1(D[5]), .A2(n1), .ZN(TMP_D[5]) );
  AND2_X1 U35 ( .A1(D[6]), .A2(n1), .ZN(TMP_D[6]) );
  AND2_X1 U36 ( .A1(D[7]), .A2(n1), .ZN(TMP_D[7]) );
  AND2_X1 U37 ( .A1(D[8]), .A2(n1), .ZN(TMP_D[8]) );
  AND2_X1 U38 ( .A1(D[31]), .A2(n1), .ZN(TMP_D[31]) );
endmodule


module FD_INJ_NB32_1 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n1, n34, n35, n36;
  wire   [31:0] TMP_D;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n36), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n36), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n36), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n36), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n36), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n36), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n36), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n36), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n35), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n35), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n35), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n35), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n35), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n35), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n35), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n35), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n35), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n35), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n35), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n35), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n34), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n34), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n34), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n34), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n34), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n34), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n34), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n34), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n34), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n34), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n34), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n34), .Q(Q[0]) );
  CLKBUF_X1 U3 ( .A(INJ_ZERO), .Z(n1) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
  BUF_X1 U6 ( .A(RESET), .Z(n36) );
  AND2_X1 U7 ( .A1(D[25]), .A2(INJ_ZERO), .ZN(TMP_D[25]) );
  AND2_X1 U8 ( .A1(D[26]), .A2(INJ_ZERO), .ZN(TMP_D[26]) );
  AND2_X1 U9 ( .A1(D[27]), .A2(INJ_ZERO), .ZN(TMP_D[27]) );
  AND2_X1 U10 ( .A1(D[28]), .A2(INJ_ZERO), .ZN(TMP_D[28]) );
  AND2_X1 U11 ( .A1(D[29]), .A2(INJ_ZERO), .ZN(TMP_D[29]) );
  AND2_X1 U12 ( .A1(D[30]), .A2(INJ_ZERO), .ZN(TMP_D[30]) );
  AND2_X1 U13 ( .A1(D[31]), .A2(n1), .ZN(TMP_D[31]) );
  AND2_X1 U14 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U15 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U16 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
  AND2_X1 U17 ( .A1(D[10]), .A2(INJ_ZERO), .ZN(TMP_D[10]) );
  AND2_X1 U18 ( .A1(D[11]), .A2(INJ_ZERO), .ZN(TMP_D[11]) );
  AND2_X1 U19 ( .A1(D[12]), .A2(INJ_ZERO), .ZN(TMP_D[12]) );
  AND2_X1 U20 ( .A1(D[13]), .A2(INJ_ZERO), .ZN(TMP_D[13]) );
  AND2_X1 U21 ( .A1(D[14]), .A2(INJ_ZERO), .ZN(TMP_D[14]) );
  AND2_X1 U22 ( .A1(D[15]), .A2(n1), .ZN(TMP_D[15]) );
  AND2_X1 U23 ( .A1(D[16]), .A2(n1), .ZN(TMP_D[16]) );
  AND2_X1 U24 ( .A1(D[17]), .A2(n1), .ZN(TMP_D[17]) );
  AND2_X1 U25 ( .A1(D[18]), .A2(n1), .ZN(TMP_D[18]) );
  AND2_X1 U26 ( .A1(D[19]), .A2(INJ_ZERO), .ZN(TMP_D[19]) );
  AND2_X1 U27 ( .A1(D[20]), .A2(INJ_ZERO), .ZN(TMP_D[20]) );
  AND2_X1 U28 ( .A1(D[21]), .A2(INJ_ZERO), .ZN(TMP_D[21]) );
  AND2_X1 U29 ( .A1(D[22]), .A2(INJ_ZERO), .ZN(TMP_D[22]) );
  AND2_X1 U30 ( .A1(D[23]), .A2(INJ_ZERO), .ZN(TMP_D[23]) );
  AND2_X1 U31 ( .A1(D[24]), .A2(INJ_ZERO), .ZN(TMP_D[24]) );
  AND2_X1 U32 ( .A1(n1), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U33 ( .A1(D[3]), .A2(n1), .ZN(TMP_D[3]) );
  AND2_X1 U34 ( .A1(D[4]), .A2(n1), .ZN(TMP_D[4]) );
  AND2_X1 U35 ( .A1(D[5]), .A2(n1), .ZN(TMP_D[5]) );
  AND2_X1 U36 ( .A1(D[6]), .A2(n1), .ZN(TMP_D[6]) );
  AND2_X1 U37 ( .A1(D[7]), .A2(n1), .ZN(TMP_D[7]) );
  AND2_X1 U38 ( .A1(D[8]), .A2(n1), .ZN(TMP_D[8]) );
endmodule


module SIGN_EXT_NB32_0 ( A, US, JMP, Y );
  input [25:0] A;
  output [31:0] Y;
  input US, JMP;
  wire   \Y[25] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  assign Y[31] = \Y[25] ;
  assign Y[30] = \Y[25] ;
  assign Y[29] = \Y[25] ;
  assign Y[28] = \Y[25] ;
  assign Y[27] = \Y[25] ;
  assign Y[26] = \Y[25] ;
  assign Y[25] = \Y[25] ;
  assign Y[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND2_X1 U2 ( .A1(n2), .A2(n12), .ZN(Y[16]) );
  NAND2_X1 U3 ( .A1(A[16]), .A2(JMP), .ZN(n12) );
  NAND2_X1 U4 ( .A1(n2), .A2(n11), .ZN(Y[17]) );
  NAND2_X1 U5 ( .A1(A[17]), .A2(JMP), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n2), .A2(n10), .ZN(Y[18]) );
  NAND2_X1 U7 ( .A1(A[18]), .A2(JMP), .ZN(n10) );
  NAND2_X1 U8 ( .A1(n2), .A2(n9), .ZN(Y[19]) );
  NAND2_X1 U9 ( .A1(A[19]), .A2(JMP), .ZN(n9) );
  NAND2_X1 U10 ( .A1(n2), .A2(n8), .ZN(Y[20]) );
  NAND2_X1 U11 ( .A1(A[20]), .A2(JMP), .ZN(n8) );
  NAND2_X1 U12 ( .A1(n2), .A2(n7), .ZN(Y[21]) );
  NAND2_X1 U13 ( .A1(A[21]), .A2(JMP), .ZN(n7) );
  NAND2_X1 U14 ( .A1(n2), .A2(n6), .ZN(Y[22]) );
  NAND2_X1 U15 ( .A1(A[22]), .A2(JMP), .ZN(n6) );
  NAND2_X1 U16 ( .A1(n2), .A2(n5), .ZN(Y[23]) );
  NAND2_X1 U17 ( .A1(A[23]), .A2(JMP), .ZN(n5) );
  NAND2_X1 U18 ( .A1(n2), .A2(n4), .ZN(Y[24]) );
  NAND2_X1 U19 ( .A1(A[24]), .A2(JMP), .ZN(n4) );
  NAND2_X1 U20 ( .A1(n13), .A2(\A[15] ), .ZN(n2) );
  NOR2_X1 U21 ( .A1(US), .A2(JMP), .ZN(n13) );
  NAND2_X1 U22 ( .A1(n2), .A2(n3), .ZN(\Y[25] ) );
  NAND2_X1 U23 ( .A1(JMP), .A2(A[25]), .ZN(n3) );
endmodule


module FD_INJ_NB32_2 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n1, n34, n35, n36, n37;
  wire   [31:0] TMP_D;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n37), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n37), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n37), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n37), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n37), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n37), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n37), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n37), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n36), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n36), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n36), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n36), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n36), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n36), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n36), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n36), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n36), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n36), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n36), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n36), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n35), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n35), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n35), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n35), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n35), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n35), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n35), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n35), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n35), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n35), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n35), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n35), .Q(Q[0]) );
  BUF_X1 U3 ( .A(RESET), .Z(n35) );
  BUF_X1 U4 ( .A(RESET), .Z(n36) );
  BUF_X1 U5 ( .A(RESET), .Z(n37) );
  BUF_X1 U6 ( .A(INJ_ZERO), .Z(n1) );
  BUF_X1 U7 ( .A(INJ_ZERO), .Z(n34) );
  AND2_X1 U8 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U9 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U10 ( .A1(D[2]), .A2(n1), .ZN(TMP_D[2]) );
  AND2_X1 U11 ( .A1(D[10]), .A2(INJ_ZERO), .ZN(TMP_D[10]) );
  AND2_X1 U12 ( .A1(D[11]), .A2(INJ_ZERO), .ZN(TMP_D[11]) );
  AND2_X1 U13 ( .A1(D[12]), .A2(INJ_ZERO), .ZN(TMP_D[12]) );
  AND2_X1 U14 ( .A1(D[13]), .A2(INJ_ZERO), .ZN(TMP_D[13]) );
  AND2_X1 U15 ( .A1(D[14]), .A2(INJ_ZERO), .ZN(TMP_D[14]) );
  AND2_X1 U16 ( .A1(D[15]), .A2(n34), .ZN(TMP_D[15]) );
  AND2_X1 U17 ( .A1(D[16]), .A2(n34), .ZN(TMP_D[16]) );
  AND2_X1 U18 ( .A1(D[17]), .A2(n34), .ZN(TMP_D[17]) );
  AND2_X1 U19 ( .A1(D[18]), .A2(n34), .ZN(TMP_D[18]) );
  AND2_X1 U20 ( .A1(D[19]), .A2(INJ_ZERO), .ZN(TMP_D[19]) );
  AND2_X1 U21 ( .A1(D[20]), .A2(n1), .ZN(TMP_D[20]) );
  AND2_X1 U22 ( .A1(D[21]), .A2(n1), .ZN(TMP_D[21]) );
  AND2_X1 U23 ( .A1(D[22]), .A2(n1), .ZN(TMP_D[22]) );
  AND2_X1 U24 ( .A1(D[23]), .A2(n1), .ZN(TMP_D[23]) );
  AND2_X1 U25 ( .A1(D[24]), .A2(n1), .ZN(TMP_D[24]) );
  AND2_X1 U26 ( .A1(D[25]), .A2(n1), .ZN(TMP_D[25]) );
  AND2_X1 U27 ( .A1(D[26]), .A2(n1), .ZN(TMP_D[26]) );
  AND2_X1 U28 ( .A1(D[27]), .A2(n1), .ZN(TMP_D[27]) );
  AND2_X1 U29 ( .A1(D[28]), .A2(n1), .ZN(TMP_D[28]) );
  AND2_X1 U30 ( .A1(D[29]), .A2(n1), .ZN(TMP_D[29]) );
  AND2_X1 U31 ( .A1(D[30]), .A2(n1), .ZN(TMP_D[30]) );
  AND2_X1 U32 ( .A1(n34), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U33 ( .A1(D[3]), .A2(n34), .ZN(TMP_D[3]) );
  AND2_X1 U34 ( .A1(D[4]), .A2(n34), .ZN(TMP_D[4]) );
  AND2_X1 U35 ( .A1(D[5]), .A2(n34), .ZN(TMP_D[5]) );
  AND2_X1 U36 ( .A1(D[6]), .A2(n34), .ZN(TMP_D[6]) );
  AND2_X1 U37 ( .A1(D[7]), .A2(n34), .ZN(TMP_D[7]) );
  AND2_X1 U38 ( .A1(D[8]), .A2(n34), .ZN(TMP_D[8]) );
  AND2_X1 U39 ( .A1(D[31]), .A2(n34), .ZN(TMP_D[31]) );
endmodule


module FD_INJ_NB32_3 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n1, n34, n35, n36, n37;
  wire   [31:0] TMP_D;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n37), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n37), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n37), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n37), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n37), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n37), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n37), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n37), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n36), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n36), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n36), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n36), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n36), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n36), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n36), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n36), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n36), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n36), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n36), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n36), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n35), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n35), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n35), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n35), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n35), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n35), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n35), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n35), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n35), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n35), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n35), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n35), .Q(Q[0]) );
  BUF_X1 U3 ( .A(RESET), .Z(n35) );
  BUF_X1 U4 ( .A(RESET), .Z(n36) );
  BUF_X1 U5 ( .A(RESET), .Z(n37) );
  AND2_X1 U6 ( .A1(D[0]), .A2(n1), .ZN(TMP_D[0]) );
  AND2_X1 U7 ( .A1(D[1]), .A2(n1), .ZN(TMP_D[1]) );
  AND2_X1 U8 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
  AND2_X1 U9 ( .A1(D[10]), .A2(n1), .ZN(TMP_D[10]) );
  AND2_X1 U10 ( .A1(D[11]), .A2(n1), .ZN(TMP_D[11]) );
  AND2_X1 U11 ( .A1(D[12]), .A2(n1), .ZN(TMP_D[12]) );
  AND2_X1 U12 ( .A1(D[13]), .A2(n1), .ZN(TMP_D[13]) );
  AND2_X1 U13 ( .A1(D[14]), .A2(n1), .ZN(TMP_D[14]) );
  AND2_X1 U14 ( .A1(D[15]), .A2(n1), .ZN(TMP_D[15]) );
  AND2_X1 U15 ( .A1(D[16]), .A2(n1), .ZN(TMP_D[16]) );
  AND2_X1 U16 ( .A1(D[17]), .A2(n1), .ZN(TMP_D[17]) );
  AND2_X1 U17 ( .A1(D[18]), .A2(n1), .ZN(TMP_D[18]) );
  AND2_X1 U18 ( .A1(D[19]), .A2(n1), .ZN(TMP_D[19]) );
  AND2_X1 U19 ( .A1(D[20]), .A2(INJ_ZERO), .ZN(TMP_D[20]) );
  AND2_X1 U20 ( .A1(D[21]), .A2(INJ_ZERO), .ZN(TMP_D[21]) );
  AND2_X1 U21 ( .A1(D[22]), .A2(INJ_ZERO), .ZN(TMP_D[22]) );
  AND2_X1 U22 ( .A1(D[23]), .A2(INJ_ZERO), .ZN(TMP_D[23]) );
  AND2_X1 U23 ( .A1(D[24]), .A2(INJ_ZERO), .ZN(TMP_D[24]) );
  AND2_X1 U24 ( .A1(D[25]), .A2(INJ_ZERO), .ZN(TMP_D[25]) );
  AND2_X1 U25 ( .A1(D[26]), .A2(n34), .ZN(TMP_D[26]) );
  AND2_X1 U26 ( .A1(D[27]), .A2(n34), .ZN(TMP_D[27]) );
  AND2_X1 U27 ( .A1(D[28]), .A2(n34), .ZN(TMP_D[28]) );
  AND2_X1 U28 ( .A1(D[29]), .A2(n34), .ZN(TMP_D[29]) );
  AND2_X1 U29 ( .A1(D[30]), .A2(INJ_ZERO), .ZN(TMP_D[30]) );
  AND2_X1 U30 ( .A1(D[6]), .A2(n34), .ZN(TMP_D[6]) );
  AND2_X1 U31 ( .A1(D[31]), .A2(n34), .ZN(TMP_D[31]) );
  AND2_X1 U32 ( .A1(D[3]), .A2(n34), .ZN(TMP_D[3]) );
  AND2_X1 U33 ( .A1(D[7]), .A2(n34), .ZN(TMP_D[7]) );
  AND2_X1 U34 ( .A1(D[4]), .A2(n34), .ZN(TMP_D[4]) );
  AND2_X1 U35 ( .A1(D[8]), .A2(n34), .ZN(TMP_D[8]) );
  AND2_X1 U36 ( .A1(D[5]), .A2(n34), .ZN(TMP_D[5]) );
  AND2_X1 U37 ( .A1(n34), .A2(D[9]), .ZN(TMP_D[9]) );
  BUF_X1 U38 ( .A(INJ_ZERO), .Z(n1) );
  BUF_X1 U39 ( .A(INJ_ZERO), .Z(n34) );
endmodule


module register_file_NB32_RS32_0 ( CLK, RESET, RD1, RD2, WR, ADD_WR, ADD_RD1, 
        ADD_RD2, DATAIN, HAZARD, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, RD1, RD2, WR;
  output HAZARD;
  wire   N4192, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297;

  DFF_X1 HAZARD_reg ( .D(N4192), .CK(CLK), .Q(HAZARD) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n3680), .CK(CLK), .Q(n3855), .QN(n274) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n3679), .CK(CLK), .Q(n3873), .QN(n281) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n3678), .CK(CLK), .Q(n3909), .QN(n295) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n3677), .CK(CLK), .Q(n3927), .QN(n302) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n3676), .CK(CLK), .Q(n3945), .QN(n309) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n3675), .CK(CLK), .Q(n3963), .QN(n316) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n3674), .CK(CLK), .Q(n3981), .QN(n323) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n3673), .CK(CLK), .Q(n3999), .QN(n330) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n3672), .CK(CLK), .Q(n4017), .QN(n337) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n3671), .CK(CLK), .Q(n4035), .QN(n344) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n3670), .CK(CLK), .Q(n4053), .QN(n351) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n3669), .CK(CLK), .Q(n4071), .QN(n358) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n3668), .CK(CLK), .Q(n4107), .QN(n372) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n3667), .CK(CLK), .Q(n4125), .QN(n379) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n3666), .CK(CLK), .Q(n4143), .QN(n386) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n3665), .CK(CLK), .Q(n4161), .QN(n393) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n3664), .CK(CLK), .Q(n4179), .QN(n400) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n3663), .CK(CLK), .Q(n4197), .QN(n407) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n3662), .CK(CLK), .Q(n4215), .QN(n414) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n3661), .CK(CLK), .Q(n4233), .QN(n421) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n3660), .CK(CLK), .Q(n4251), .QN(n428) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n3659), .CK(CLK), .Q(n4269), .QN(n435) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n3658), .CK(CLK), .Q(n3729), .QN(n225) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n3657), .CK(CLK), .Q(n3747), .QN(n232) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n3656), .CK(CLK), .Q(n3765), .QN(n239) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n3655), .CK(CLK), .Q(n3783), .QN(n246) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n3654), .CK(CLK), .Q(n3801), .QN(n253) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n3653), .CK(CLK), .Q(n3819), .QN(n260) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n3652), .CK(CLK), .Q(n3837), .QN(n267) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n3651), .CK(CLK), .Q(n3891), .QN(n288) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n3650), .CK(CLK), .Q(n4089), .QN(n365) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n3649), .CK(CLK), .Q(n4287), .QN(n442) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n3648), .CK(CLK), .Q(n3854), .QN(n50) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n3647), .CK(CLK), .Q(n3872), .QN(n57) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n3646), .CK(CLK), .Q(n3908), .QN(n71) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n3645), .CK(CLK), .Q(n3926), .QN(n78) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n3644), .CK(CLK), .Q(n3944), .QN(n85) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n3643), .CK(CLK), .Q(n3962), .QN(n92) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n3642), .CK(CLK), .Q(n3980), .QN(n99) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n3641), .CK(CLK), .Q(n3998), .QN(n106) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n3640), .CK(CLK), .Q(n4016), .QN(n113) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n3639), .CK(CLK), .Q(n4034), .QN(n120) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n3638), .CK(CLK), .Q(n4052), .QN(n127) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n3637), .CK(CLK), .Q(n4070), .QN(n134) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n3636), .CK(CLK), .Q(n4106), .QN(n148) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n3635), .CK(CLK), .Q(n4124), .QN(n155) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n3634), .CK(CLK), .Q(n4142), .QN(n162) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n3633), .CK(CLK), .Q(n4160), .QN(n169) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n3632), .CK(CLK), .Q(n4178), .QN(n176) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n3631), .CK(CLK), .Q(n4196), .QN(n183) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n3630), .CK(CLK), .Q(n4214), .QN(n190) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n3629), .CK(CLK), .Q(n4232), .QN(n197) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n3628), .CK(CLK), .Q(n4250), .QN(n204) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n3627), .CK(CLK), .Q(n4268), .QN(n211) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n3626), .CK(CLK), .Q(n3728), .QN(n1) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n3625), .CK(CLK), .Q(n3746), .QN(n8) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n3624), .CK(CLK), .Q(n3764), .QN(n15) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n3623), .CK(CLK), .Q(n3782), .QN(n22) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n3622), .CK(CLK), .Q(n3800), .QN(n29) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n3621), .CK(CLK), .Q(n3818), .QN(n36) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n3620), .CK(CLK), .Q(n3836), .QN(n43) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n3619), .CK(CLK), .Q(n3890), .QN(n64) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n3618), .CK(CLK), .Q(n4088), .QN(n141) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n3617), .CK(CLK), .Q(n4286), .QN(n218) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n3616), .CK(CLK), .Q(n873) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n3615), .CK(CLK), .Q(n875) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n3614), .CK(CLK), .Q(n876) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n3613), .CK(CLK), .Q(n877) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n3612), .CK(CLK), .Q(n878) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n3611), .CK(CLK), .Q(n879) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n3610), .CK(CLK), .Q(n880) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n3609), .CK(CLK), .Q(n881) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n3608), .CK(CLK), .Q(n882) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n3607), .CK(CLK), .Q(n883) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n3606), .CK(CLK), .Q(n884) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n3605), .CK(CLK), .Q(n885) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n3604), .CK(CLK), .Q(n886) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n3603), .CK(CLK), .Q(n887) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n3602), .CK(CLK), .Q(n888) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n3601), .CK(CLK), .Q(n889) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n3600), .CK(CLK), .Q(n890) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n3599), .CK(CLK), .Q(n891) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n3598), .CK(CLK), .Q(n892) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n3597), .CK(CLK), .Q(n893) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n3596), .CK(CLK), .Q(n894) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n3595), .CK(CLK), .Q(n895) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n3594), .CK(CLK), .Q(n896) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n3593), .CK(CLK), .Q(n897) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n3592), .CK(CLK), .Q(n898) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n3591), .CK(CLK), .Q(n899) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n3590), .CK(CLK), .Q(n900) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n3589), .CK(CLK), .Q(n901) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n3588), .CK(CLK), .Q(n902) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n3587), .CK(CLK), .Q(n903) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n3586), .CK(CLK), .Q(n904) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n3585), .CK(CLK), .Q(n905) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n3584), .CK(CLK), .Q(n907) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n3583), .CK(CLK), .Q(n909) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n3582), .CK(CLK), .Q(n910) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n3581), .CK(CLK), .Q(n911) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n3580), .CK(CLK), .Q(n912) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n3579), .CK(CLK), .Q(n913) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n3578), .CK(CLK), .Q(n914) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n3577), .CK(CLK), .Q(n915) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n3576), .CK(CLK), .Q(n916) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n3575), .CK(CLK), .Q(n917) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n3574), .CK(CLK), .Q(n918) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n3573), .CK(CLK), .Q(n919) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n3572), .CK(CLK), .Q(n920) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n3571), .CK(CLK), .Q(n921) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n3570), .CK(CLK), .Q(n922) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n3569), .CK(CLK), .Q(n923) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n3568), .CK(CLK), .Q(n924) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n3567), .CK(CLK), .Q(n925) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n3566), .CK(CLK), .Q(n926) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n3565), .CK(CLK), .Q(n927) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n3564), .CK(CLK), .Q(n928) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n3563), .CK(CLK), .Q(n929) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n3562), .CK(CLK), .Q(n930) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n3561), .CK(CLK), .Q(n931) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n3560), .CK(CLK), .Q(n932) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n3559), .CK(CLK), .Q(n933) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n3558), .CK(CLK), .Q(n934) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n3557), .CK(CLK), .Q(n935) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n3556), .CK(CLK), .Q(n936) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n3555), .CK(CLK), .Q(n937) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n3554), .CK(CLK), .Q(n938) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n3553), .CK(CLK), .Q(n939) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n3552), .CK(CLK), .Q(n3853), .QN(n275) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n3551), .CK(CLK), .Q(n3871), .QN(n282) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n3550), .CK(CLK), .Q(n3907), .QN(n296) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n3549), .CK(CLK), .Q(n3925), .QN(n303) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n3548), .CK(CLK), .Q(n3943), .QN(n310) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n3547), .CK(CLK), .Q(n3961), .QN(n317) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n3546), .CK(CLK), .Q(n3979), .QN(n324) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n3545), .CK(CLK), .Q(n3997), .QN(n331) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n3544), .CK(CLK), .Q(n4015), .QN(n338) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n3543), .CK(CLK), .Q(n4033), .QN(n345) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n3542), .CK(CLK), .Q(n4051), .QN(n352) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n3541), .CK(CLK), .Q(n4069), .QN(n359) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n3540), .CK(CLK), .Q(n4105), .QN(n373) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n3539), .CK(CLK), .Q(n4123), .QN(n380) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n3538), .CK(CLK), .Q(n4141), .QN(n387) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n3537), .CK(CLK), .Q(n4159), .QN(n394) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n3536), .CK(CLK), .Q(n4177), .QN(n401) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n3535), .CK(CLK), .Q(n4195), .QN(n408) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n3534), .CK(CLK), .Q(n4213), .QN(n415) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n3533), .CK(CLK), .Q(n4231), .QN(n422) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n3532), .CK(CLK), .Q(n4249), .QN(n429) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n3531), .CK(CLK), .Q(n4267), .QN(n436) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n3530), .CK(CLK), .Q(n3727), .QN(n226) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n3529), .CK(CLK), .Q(n3745), .QN(n233) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n3528), .CK(CLK), .Q(n3763), .QN(n240) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n3527), .CK(CLK), .Q(n3781), .QN(n247) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n3526), .CK(CLK), .Q(n3799), .QN(n254) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n3525), .CK(CLK), .Q(n3817), .QN(n261) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n3524), .CK(CLK), .Q(n3835), .QN(n268) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n3523), .CK(CLK), .Q(n3889), .QN(n289) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n3522), .CK(CLK), .Q(n4087), .QN(n366) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n3521), .CK(CLK), .Q(n4285), .QN(n443) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n3520), .CK(CLK), .Q(n3852), .QN(n51) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n3519), .CK(CLK), .Q(n3870), .QN(n58) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n3518), .CK(CLK), .Q(n3906), .QN(n72) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n3517), .CK(CLK), .Q(n3924), .QN(n79) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n3516), .CK(CLK), .Q(n3942), .QN(n86) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n3515), .CK(CLK), .Q(n3960), .QN(n93) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n3514), .CK(CLK), .Q(n3978), .QN(n100) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n3513), .CK(CLK), .Q(n3996), .QN(n107) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n3512), .CK(CLK), .Q(n4014), .QN(n114) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n3511), .CK(CLK), .Q(n4032), .QN(n121) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n3510), .CK(CLK), .Q(n4050), .QN(n128) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n3509), .CK(CLK), .Q(n4068), .QN(n135) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n3508), .CK(CLK), .Q(n4104), .QN(n149) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n3507), .CK(CLK), .Q(n4122), .QN(n156) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n3506), .CK(CLK), .Q(n4140), .QN(n163) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n3505), .CK(CLK), .Q(n4158), .QN(n170) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n3504), .CK(CLK), .Q(n4176), .QN(n177) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n3503), .CK(CLK), .Q(n4194), .QN(n184) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n3502), .CK(CLK), .Q(n4212), .QN(n191) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n3501), .CK(CLK), .Q(n4230), .QN(n198) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n3500), .CK(CLK), .Q(n4248), .QN(n205) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n3499), .CK(CLK), .Q(n4266), .QN(n212) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n3498), .CK(CLK), .Q(n3726), .QN(n2) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n3497), .CK(CLK), .Q(n3744), .QN(n9) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n3496), .CK(CLK), .Q(n3762), .QN(n16) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n3495), .CK(CLK), .Q(n3780), .QN(n23) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n3494), .CK(CLK), .Q(n3798), .QN(n30) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n3493), .CK(CLK), .Q(n3816), .QN(n37) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n3492), .CK(CLK), .Q(n3834), .QN(n44) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n3491), .CK(CLK), .Q(n3888), .QN(n65) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n3490), .CK(CLK), .Q(n4086), .QN(n142) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n3489), .CK(CLK), .Q(n4284), .QN(n219) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n3488), .CK(CLK), .Q(n947) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n3487), .CK(CLK), .Q(n949) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n3486), .CK(CLK), .Q(n950) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n3485), .CK(CLK), .Q(n951) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n3484), .CK(CLK), .Q(n952) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n3483), .CK(CLK), .Q(n953) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n3482), .CK(CLK), .Q(n954) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n3481), .CK(CLK), .Q(n955) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n3480), .CK(CLK), .Q(n956) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n3479), .CK(CLK), .Q(n957) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n3478), .CK(CLK), .Q(n958) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n3477), .CK(CLK), .Q(n959) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n3476), .CK(CLK), .Q(n960) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n3475), .CK(CLK), .Q(n961) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n3474), .CK(CLK), .Q(n962) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n3473), .CK(CLK), .Q(n963) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n3472), .CK(CLK), .Q(n964) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n3471), .CK(CLK), .Q(n965) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n3470), .CK(CLK), .Q(n966) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n3469), .CK(CLK), .Q(n967) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n3468), .CK(CLK), .Q(n968) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n3467), .CK(CLK), .Q(n969) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n3466), .CK(CLK), .Q(n970) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n3465), .CK(CLK), .Q(n971) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n3464), .CK(CLK), .Q(n972) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n3463), .CK(CLK), .Q(n973) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n3462), .CK(CLK), .Q(n974) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n3461), .CK(CLK), .Q(n975) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n3460), .CK(CLK), .Q(n976) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n3459), .CK(CLK), .Q(n977) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n3458), .CK(CLK), .Q(n978) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n3457), .CK(CLK), .Q(n979) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n3456), .CK(CLK), .Q(n980) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n3455), .CK(CLK), .Q(n982) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n3454), .CK(CLK), .Q(n983) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n3453), .CK(CLK), .Q(n984) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n3452), .CK(CLK), .Q(n985) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n3451), .CK(CLK), .Q(n986) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n3450), .CK(CLK), .Q(n987) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n3449), .CK(CLK), .Q(n988) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n3448), .CK(CLK), .Q(n989) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n3447), .CK(CLK), .Q(n990) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n3446), .CK(CLK), .Q(n991) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n3445), .CK(CLK), .Q(n992) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n3444), .CK(CLK), .Q(n993) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n3443), .CK(CLK), .Q(n994) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n3442), .CK(CLK), .Q(n995) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n3441), .CK(CLK), .Q(n996) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n3440), .CK(CLK), .Q(n997) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n3439), .CK(CLK), .Q(n998) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n3438), .CK(CLK), .Q(n999) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n3437), .CK(CLK), .Q(n1000) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n3436), .CK(CLK), .Q(n1001) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n3435), .CK(CLK), .Q(n1002) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n3434), .CK(CLK), .Q(n1003) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n3433), .CK(CLK), .Q(n1004) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n3432), .CK(CLK), .Q(n1005) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n3431), .CK(CLK), .Q(n1006) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n3430), .CK(CLK), .Q(n1007) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n3429), .CK(CLK), .Q(n1008) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n3428), .CK(CLK), .Q(n1009) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n3427), .CK(CLK), .Q(n1010) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n3426), .CK(CLK), .Q(n1011) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n3425), .CK(CLK), .Q(n1012) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n3424), .CK(CLK), .Q(n3851), .QN(n276) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n3423), .CK(CLK), .Q(n3869), .QN(n283) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n3422), .CK(CLK), .Q(n3905), .QN(n297) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n3421), .CK(CLK), .Q(n3923), .QN(n304) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n3420), .CK(CLK), .Q(n3941), .QN(n311) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n3419), .CK(CLK), .Q(n3959), .QN(n318) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n3418), .CK(CLK), .Q(n3977), .QN(n325) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n3417), .CK(CLK), .Q(n3995), .QN(n332) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n3416), .CK(CLK), .Q(n4013), .QN(n339) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n3415), .CK(CLK), .Q(n4031), .QN(n346) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n3414), .CK(CLK), .Q(n4049), .QN(n353) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n3413), .CK(CLK), .Q(n4067), .QN(n360) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n3412), .CK(CLK), .Q(n4103), .QN(n374) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n3411), .CK(CLK), .Q(n4121), .QN(n381) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n3410), .CK(CLK), .Q(n4139), .QN(n388) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n3409), .CK(CLK), .Q(n4157), .QN(n395) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n3408), .CK(CLK), .Q(n4175), .QN(n402) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n3407), .CK(CLK), .Q(n4193), .QN(n409) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n3406), .CK(CLK), .Q(n4211), .QN(n416) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n3405), .CK(CLK), .Q(n4229), .QN(n423) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n3404), .CK(CLK), .Q(n4247), .QN(n430) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n3403), .CK(CLK), .Q(n4265), .QN(n437) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n3402), .CK(CLK), .Q(n3725), .QN(n227) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n3401), .CK(CLK), .Q(n3743), .QN(n234) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n3400), .CK(CLK), .Q(n3761), .QN(n241) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n3399), .CK(CLK), .Q(n3779), .QN(n248) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n3398), .CK(CLK), .Q(n3797), .QN(n255) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n3397), .CK(CLK), .Q(n3815), .QN(n262) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n3396), .CK(CLK), .Q(n3833), .QN(n269) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n3395), .CK(CLK), .Q(n3887), .QN(n290) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n3394), .CK(CLK), .Q(n4085), .QN(n367) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n3393), .CK(CLK), .Q(n4283), .QN(n444) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n3392), .CK(CLK), .Q(n3850), .QN(n52) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n3391), .CK(CLK), .Q(n3868), .QN(n59) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n3390), .CK(CLK), .Q(n3904), .QN(n73) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n3389), .CK(CLK), .Q(n3922), .QN(n80) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n3388), .CK(CLK), .Q(n3940), .QN(n87) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n3387), .CK(CLK), .Q(n3958), .QN(n94) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n3386), .CK(CLK), .Q(n3976), .QN(n101) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n3385), .CK(CLK), .Q(n3994), .QN(n108) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n3384), .CK(CLK), .Q(n4012), .QN(n115) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n3383), .CK(CLK), .Q(n4030), .QN(n122) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n3382), .CK(CLK), .Q(n4048), .QN(n129) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n3381), .CK(CLK), .Q(n4066), .QN(n136) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n3380), .CK(CLK), .Q(n4102), .QN(n150) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n3379), .CK(CLK), .Q(n4120), .QN(n157) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n3378), .CK(CLK), .Q(n4138), .QN(n164) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n3377), .CK(CLK), .Q(n4156), .QN(n171) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n3376), .CK(CLK), .Q(n4174), .QN(n178) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n3375), .CK(CLK), .Q(n4192), .QN(n185) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n3374), .CK(CLK), .Q(n4210), .QN(n192) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n3373), .CK(CLK), .Q(n4228), .QN(n199) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n3372), .CK(CLK), .Q(n4246), .QN(n206) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n3371), .CK(CLK), .Q(n4264), .QN(n213) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n3370), .CK(CLK), .Q(n3724), .QN(n3) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n3369), .CK(CLK), .Q(n3742), .QN(n10) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n3368), .CK(CLK), .Q(n3760), .QN(n17) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n3367), .CK(CLK), .Q(n3778), .QN(n24) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n3366), .CK(CLK), .Q(n3796), .QN(n31) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n3365), .CK(CLK), .Q(n3814), .QN(n38) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n3364), .CK(CLK), .Q(n3832), .QN(n45) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n3363), .CK(CLK), .Q(n3886), .QN(n66) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n3362), .CK(CLK), .Q(n4084), .QN(n143) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n3361), .CK(CLK), .Q(n4282), .QN(n220) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n3360), .CK(CLK), .Q(n1016) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n3359), .CK(CLK), .Q(n1018) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n3358), .CK(CLK), .Q(n1019) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n3357), .CK(CLK), .Q(n1020) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n3356), .CK(CLK), .Q(n1021) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n3355), .CK(CLK), .Q(n1022) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n3354), .CK(CLK), .Q(n1023) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n3353), .CK(CLK), .Q(n1024) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n3352), .CK(CLK), .Q(n1025) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n3351), .CK(CLK), .Q(n1026) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n3350), .CK(CLK), .Q(n1027) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n3349), .CK(CLK), .Q(n1028) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n3348), .CK(CLK), .Q(n1029) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n3347), .CK(CLK), .Q(n1030) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n3346), .CK(CLK), .Q(n1031) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n3345), .CK(CLK), .Q(n1032) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n3344), .CK(CLK), .Q(n1033) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n3343), .CK(CLK), .Q(n1034) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n3342), .CK(CLK), .Q(n1035) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n3341), .CK(CLK), .Q(n1036) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n3340), .CK(CLK), .Q(n1037) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n3339), .CK(CLK), .Q(n1038) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n3338), .CK(CLK), .Q(n1039) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n3337), .CK(CLK), .Q(n1040) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n3336), .CK(CLK), .Q(n1041) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n3335), .CK(CLK), .Q(n1042) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n3334), .CK(CLK), .Q(n1043) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n3333), .CK(CLK), .Q(n1044) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n3332), .CK(CLK), .Q(n1045) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n3331), .CK(CLK), .Q(n1046) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n3330), .CK(CLK), .Q(n1047) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n3329), .CK(CLK), .Q(n1048) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n3328), .CK(CLK), .Q(n1049) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n3327), .CK(CLK), .Q(n1051) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n3326), .CK(CLK), .Q(n1052) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n3325), .CK(CLK), .Q(n1053) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n3324), .CK(CLK), .Q(n1054) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n3323), .CK(CLK), .Q(n1055) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n3322), .CK(CLK), .Q(n1056) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n3321), .CK(CLK), .Q(n1057) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n3320), .CK(CLK), .Q(n1058) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n3319), .CK(CLK), .Q(n1059) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n3318), .CK(CLK), .Q(n1060) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n3317), .CK(CLK), .Q(n1061) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n3316), .CK(CLK), .Q(n1062) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n3315), .CK(CLK), .Q(n1063) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n3314), .CK(CLK), .Q(n1064) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n3313), .CK(CLK), .Q(n1065) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n3312), .CK(CLK), .Q(n1066) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n3311), .CK(CLK), .Q(n1067) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n3310), .CK(CLK), .Q(n1068) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n3309), .CK(CLK), .Q(n1069) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n3308), .CK(CLK), .Q(n1070) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n3307), .CK(CLK), .Q(n1071) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n3306), .CK(CLK), .Q(n1072) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n3305), .CK(CLK), .Q(n1073) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n3304), .CK(CLK), .Q(n1074) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n3303), .CK(CLK), .Q(n1075) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n3302), .CK(CLK), .Q(n1076) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n3301), .CK(CLK), .Q(n1077) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n3300), .CK(CLK), .Q(n1078) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n3299), .CK(CLK), .Q(n1079) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n3298), .CK(CLK), .Q(n1080) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n3297), .CK(CLK), .Q(n1081) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n3296), .CK(CLK), .Q(n3849), .QN(n277)
         );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n3295), .CK(CLK), .Q(n3867), .QN(n284)
         );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n3294), .CK(CLK), .Q(n3903), .QN(n298)
         );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n3293), .CK(CLK), .Q(n3921), .QN(n305)
         );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n3292), .CK(CLK), .Q(n3939), .QN(n312)
         );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n3291), .CK(CLK), .Q(n3957), .QN(n319)
         );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n3290), .CK(CLK), .Q(n3975), .QN(n326)
         );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n3289), .CK(CLK), .Q(n3993), .QN(n333)
         );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n3288), .CK(CLK), .Q(n4011), .QN(n340)
         );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n3287), .CK(CLK), .Q(n4029), .QN(n347)
         );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n3286), .CK(CLK), .Q(n4047), .QN(n354)
         );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n3285), .CK(CLK), .Q(n4065), .QN(n361)
         );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n3284), .CK(CLK), .Q(n4101), .QN(n375)
         );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n3283), .CK(CLK), .Q(n4119), .QN(n382)
         );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n3282), .CK(CLK), .Q(n4137), .QN(n389)
         );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n3281), .CK(CLK), .Q(n4155), .QN(n396)
         );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n3280), .CK(CLK), .Q(n4173), .QN(n403)
         );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n3279), .CK(CLK), .Q(n4191), .QN(n410)
         );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n3278), .CK(CLK), .Q(n4209), .QN(n417)
         );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n3277), .CK(CLK), .Q(n4227), .QN(n424)
         );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n3276), .CK(CLK), .Q(n4245), .QN(n431)
         );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n3275), .CK(CLK), .Q(n4263), .QN(n438)
         );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n3274), .CK(CLK), .Q(n3723), .QN(n228) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n3273), .CK(CLK), .Q(n3741), .QN(n235) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n3272), .CK(CLK), .Q(n3759), .QN(n242) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n3271), .CK(CLK), .Q(n3777), .QN(n249) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n3270), .CK(CLK), .Q(n3795), .QN(n256) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n3269), .CK(CLK), .Q(n3813), .QN(n263) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n3268), .CK(CLK), .Q(n3831), .QN(n270) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n3267), .CK(CLK), .Q(n3885), .QN(n291) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n3266), .CK(CLK), .Q(n4083), .QN(n368) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n3265), .CK(CLK), .Q(n4281), .QN(n445) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n3264), .CK(CLK), .Q(n3848), .QN(n53) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n3263), .CK(CLK), .Q(n3866), .QN(n60) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n3262), .CK(CLK), .Q(n3902), .QN(n74) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n3261), .CK(CLK), .Q(n3920), .QN(n81) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n3260), .CK(CLK), .Q(n3938), .QN(n88) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n3259), .CK(CLK), .Q(n3956), .QN(n95) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n3258), .CK(CLK), .Q(n3974), .QN(n102)
         );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n3257), .CK(CLK), .Q(n3992), .QN(n109)
         );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n3256), .CK(CLK), .Q(n4010), .QN(n116)
         );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n3255), .CK(CLK), .Q(n4028), .QN(n123)
         );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n3254), .CK(CLK), .Q(n4046), .QN(n130)
         );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n3253), .CK(CLK), .Q(n4064), .QN(n137)
         );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n3252), .CK(CLK), .Q(n4100), .QN(n151)
         );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n3251), .CK(CLK), .Q(n4118), .QN(n158)
         );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n3250), .CK(CLK), .Q(n4136), .QN(n165)
         );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n3249), .CK(CLK), .Q(n4154), .QN(n172)
         );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n3248), .CK(CLK), .Q(n4172), .QN(n179)
         );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n3247), .CK(CLK), .Q(n4190), .QN(n186)
         );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n3246), .CK(CLK), .Q(n4208), .QN(n193)
         );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n3245), .CK(CLK), .Q(n4226), .QN(n200)
         );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n3244), .CK(CLK), .Q(n4244), .QN(n207)
         );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n3243), .CK(CLK), .Q(n4262), .QN(n214)
         );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n3242), .CK(CLK), .Q(n3722), .QN(n4) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n3241), .CK(CLK), .Q(n3740), .QN(n11) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n3240), .CK(CLK), .Q(n3758), .QN(n18) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n3239), .CK(CLK), .Q(n3776), .QN(n25) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n3238), .CK(CLK), .Q(n3794), .QN(n32) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n3237), .CK(CLK), .Q(n3812), .QN(n39) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n3236), .CK(CLK), .Q(n3830), .QN(n46) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n3235), .CK(CLK), .Q(n3884), .QN(n67) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n3234), .CK(CLK), .Q(n4082), .QN(n144) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n3233), .CK(CLK), .Q(n4280), .QN(n221) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n3232), .CK(CLK), .Q(n1085) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n3231), .CK(CLK), .Q(n1087) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n3230), .CK(CLK), .Q(n1088) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n3229), .CK(CLK), .Q(n1089) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n3228), .CK(CLK), .Q(n1090) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n3227), .CK(CLK), .Q(n1091) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n3226), .CK(CLK), .Q(n1092) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n3225), .CK(CLK), .Q(n1093) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n3224), .CK(CLK), .Q(n1094) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n3223), .CK(CLK), .Q(n1095) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n3222), .CK(CLK), .Q(n1096) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n3221), .CK(CLK), .Q(n1097) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n3220), .CK(CLK), .Q(n1098) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n3219), .CK(CLK), .Q(n1099) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n3218), .CK(CLK), .Q(n1100) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n3217), .CK(CLK), .Q(n1101) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n3216), .CK(CLK), .Q(n1102) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n3215), .CK(CLK), .Q(n1103) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n3214), .CK(CLK), .Q(n1104) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n3213), .CK(CLK), .Q(n1105) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n3212), .CK(CLK), .Q(n1106) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n3211), .CK(CLK), .Q(n1107) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n3210), .CK(CLK), .Q(n1108) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n3209), .CK(CLK), .Q(n1109) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n3208), .CK(CLK), .Q(n1110) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n3207), .CK(CLK), .Q(n1111) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n3206), .CK(CLK), .Q(n1112) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n3205), .CK(CLK), .Q(n1113) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n3204), .CK(CLK), .Q(n1114) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n3203), .CK(CLK), .Q(n1115) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n3202), .CK(CLK), .Q(n1116) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n3201), .CK(CLK), .Q(n1117) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n3200), .CK(CLK), .Q(n1118) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n3199), .CK(CLK), .Q(n1120) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n3198), .CK(CLK), .Q(n1121) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n3197), .CK(CLK), .Q(n1122) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n3196), .CK(CLK), .Q(n1123) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n3195), .CK(CLK), .Q(n1124) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n3194), .CK(CLK), .Q(n1125) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n3193), .CK(CLK), .Q(n1126) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n3192), .CK(CLK), .Q(n1127) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n3191), .CK(CLK), .Q(n1128) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n3190), .CK(CLK), .Q(n1129) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n3189), .CK(CLK), .Q(n1130) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n3188), .CK(CLK), .Q(n1131) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n3187), .CK(CLK), .Q(n1132) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n3186), .CK(CLK), .Q(n1133) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n3185), .CK(CLK), .Q(n1134) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n3184), .CK(CLK), .Q(n1135) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n3183), .CK(CLK), .Q(n1136) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n3182), .CK(CLK), .Q(n1137) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n3181), .CK(CLK), .Q(n1138) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n3180), .CK(CLK), .Q(n1139) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n3179), .CK(CLK), .Q(n1140) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n3178), .CK(CLK), .Q(n1141) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n3177), .CK(CLK), .Q(n1142) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n3176), .CK(CLK), .Q(n1143) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n3175), .CK(CLK), .Q(n1144) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n3174), .CK(CLK), .Q(n1145) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n3173), .CK(CLK), .Q(n1146) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n3172), .CK(CLK), .Q(n1147) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n3171), .CK(CLK), .Q(n1148) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n3170), .CK(CLK), .Q(n1149) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n3169), .CK(CLK), .Q(n1150) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n3168), .CK(CLK), .Q(n3858), .QN(n55) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n3167), .CK(CLK), .Q(n3876), .QN(n62) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n3166), .CK(CLK), .Q(n3912), .QN(n76) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n3165), .CK(CLK), .Q(n3930), .QN(n83) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n3164), .CK(CLK), .Q(n3948), .QN(n90) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n3163), .CK(CLK), .Q(n3966), .QN(n97) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n3162), .CK(CLK), .Q(n3984), .QN(n104)
         );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n3161), .CK(CLK), .Q(n4002), .QN(n111)
         );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n3160), .CK(CLK), .Q(n4020), .QN(n118)
         );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n3159), .CK(CLK), .Q(n4038), .QN(n125)
         );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n3158), .CK(CLK), .Q(n4056), .QN(n132)
         );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n3157), .CK(CLK), .Q(n4074), .QN(n139)
         );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n3156), .CK(CLK), .Q(n4110), .QN(n153)
         );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n3155), .CK(CLK), .Q(n4128), .QN(n160)
         );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n3154), .CK(CLK), .Q(n4146), .QN(n167)
         );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n3153), .CK(CLK), .Q(n4164), .QN(n174)
         );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n3152), .CK(CLK), .Q(n4182), .QN(n181)
         );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n3151), .CK(CLK), .Q(n4200), .QN(n188)
         );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n3150), .CK(CLK), .Q(n4218), .QN(n195)
         );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n3149), .CK(CLK), .Q(n4236), .QN(n202)
         );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n3148), .CK(CLK), .Q(n4254), .QN(n209)
         );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n3147), .CK(CLK), .Q(n4272), .QN(n216)
         );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n3146), .CK(CLK), .Q(n3732), .QN(n6) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n3145), .CK(CLK), .Q(n3750), .QN(n13) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n3144), .CK(CLK), .Q(n3768), .QN(n20) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n3143), .CK(CLK), .Q(n3786), .QN(n27) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n3142), .CK(CLK), .Q(n3804), .QN(n34) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n3141), .CK(CLK), .Q(n3822), .QN(n41) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n3140), .CK(CLK), .Q(n3840), .QN(n48) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n3139), .CK(CLK), .Q(n3894), .QN(n69) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n3138), .CK(CLK), .Q(n4092), .QN(n146) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n3137), .CK(CLK), .Q(n4290), .QN(n223) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n3136), .CK(CLK), .Q(n3859), .QN(n279)
         );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n3135), .CK(CLK), .Q(n3877), .QN(n286)
         );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n3134), .CK(CLK), .Q(n3913), .QN(n300)
         );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n3133), .CK(CLK), .Q(n3931), .QN(n307)
         );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n3132), .CK(CLK), .Q(n3949), .QN(n314)
         );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n3131), .CK(CLK), .Q(n3967), .QN(n321)
         );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n3130), .CK(CLK), .Q(n3985), .QN(n328)
         );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n3129), .CK(CLK), .Q(n4003), .QN(n335)
         );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n3128), .CK(CLK), .Q(n4021), .QN(n342)
         );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n3127), .CK(CLK), .Q(n4039), .QN(n349)
         );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n3126), .CK(CLK), .Q(n4057), .QN(n356)
         );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n3125), .CK(CLK), .Q(n4075), .QN(n363)
         );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n3124), .CK(CLK), .Q(n4111), .QN(n377)
         );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n3123), .CK(CLK), .Q(n4129), .QN(n384)
         );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n3122), .CK(CLK), .Q(n4147), .QN(n391)
         );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n3121), .CK(CLK), .Q(n4165), .QN(n398)
         );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n3120), .CK(CLK), .Q(n4183), .QN(n405)
         );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n3119), .CK(CLK), .Q(n4201), .QN(n412)
         );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n3118), .CK(CLK), .Q(n4219), .QN(n419)
         );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n3117), .CK(CLK), .Q(n4237), .QN(n426)
         );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n3116), .CK(CLK), .Q(n4255), .QN(n433)
         );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n3115), .CK(CLK), .Q(n4273), .QN(n440)
         );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n3114), .CK(CLK), .Q(n3733), .QN(n230) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n3113), .CK(CLK), .Q(n3751), .QN(n237) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n3112), .CK(CLK), .Q(n3769), .QN(n244) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n3111), .CK(CLK), .Q(n3787), .QN(n251) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n3110), .CK(CLK), .Q(n3805), .QN(n258) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n3109), .CK(CLK), .Q(n3823), .QN(n265) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n3108), .CK(CLK), .Q(n3841), .QN(n272) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n3107), .CK(CLK), .Q(n3895), .QN(n293) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n3106), .CK(CLK), .Q(n4093), .QN(n370) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n3105), .CK(CLK), .Q(n4291), .QN(n447) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n3104), .CK(CLK), .Q(n1155) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n3103), .CK(CLK), .Q(n1157) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n3102), .CK(CLK), .Q(n1158) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n3101), .CK(CLK), .Q(n1159) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n3100), .CK(CLK), .Q(n1160) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n3099), .CK(CLK), .Q(n1161) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n3098), .CK(CLK), .Q(n1162) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n3097), .CK(CLK), .Q(n1163) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n3096), .CK(CLK), .Q(n1164) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n3095), .CK(CLK), .Q(n1165) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n3094), .CK(CLK), .Q(n1166) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n3093), .CK(CLK), .Q(n1167) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n3092), .CK(CLK), .Q(n1168) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n3091), .CK(CLK), .Q(n1169) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n3090), .CK(CLK), .Q(n1170) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n3089), .CK(CLK), .Q(n1171) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n3088), .CK(CLK), .Q(n1172) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n3087), .CK(CLK), .Q(n1173) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n3086), .CK(CLK), .Q(n1174) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n3085), .CK(CLK), .Q(n1175) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n3084), .CK(CLK), .Q(n1176) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n3083), .CK(CLK), .Q(n1177) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n3082), .CK(CLK), .Q(n1178) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n3081), .CK(CLK), .Q(n1179) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n3080), .CK(CLK), .Q(n1180) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n3079), .CK(CLK), .Q(n1181) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n3078), .CK(CLK), .Q(n1182) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n3077), .CK(CLK), .Q(n1183) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n3076), .CK(CLK), .Q(n1184) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n3075), .CK(CLK), .Q(n1185) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n3074), .CK(CLK), .Q(n1186) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n3073), .CK(CLK), .Q(n1187) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n3072), .CK(CLK), .Q(n1188) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n3071), .CK(CLK), .Q(n1190) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n3070), .CK(CLK), .Q(n1191) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n3069), .CK(CLK), .Q(n1192) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n3068), .CK(CLK), .Q(n1193) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n3067), .CK(CLK), .Q(n1194) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n3066), .CK(CLK), .Q(n1195) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n3065), .CK(CLK), .Q(n1196) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n3064), .CK(CLK), .Q(n1197) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n3063), .CK(CLK), .Q(n1198) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n3062), .CK(CLK), .Q(n1199) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n3061), .CK(CLK), .Q(n1200) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n3060), .CK(CLK), .Q(n1201) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n3059), .CK(CLK), .Q(n1202) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n3058), .CK(CLK), .Q(n1203) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n3057), .CK(CLK), .Q(n1204) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n3056), .CK(CLK), .Q(n1205) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n3055), .CK(CLK), .Q(n1206) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n3054), .CK(CLK), .Q(n1207) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n3053), .CK(CLK), .Q(n1208) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n3052), .CK(CLK), .Q(n1209) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n3051), .CK(CLK), .Q(n1210) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n3050), .CK(CLK), .Q(n1211) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n3049), .CK(CLK), .Q(n1212) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n3048), .CK(CLK), .Q(n1213) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n3047), .CK(CLK), .Q(n1214) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n3046), .CK(CLK), .Q(n1215) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n3045), .CK(CLK), .Q(n1216) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n3044), .CK(CLK), .Q(n1217) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n3043), .CK(CLK), .Q(n1218) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n3042), .CK(CLK), .Q(n1219) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n3041), .CK(CLK), .Q(n1220) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n3040), .CK(CLK), .Q(n3856), .QN(n56) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n3039), .CK(CLK), .Q(n3874), .QN(n63) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n3038), .CK(CLK), .Q(n3910), .QN(n77) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n3037), .CK(CLK), .Q(n3928), .QN(n84) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n3036), .CK(CLK), .Q(n3946), .QN(n91) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n3035), .CK(CLK), .Q(n3964), .QN(n98) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n3034), .CK(CLK), .Q(n3982), .QN(n105)
         );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n3033), .CK(CLK), .Q(n4000), .QN(n112)
         );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n3032), .CK(CLK), .Q(n4018), .QN(n119)
         );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n3031), .CK(CLK), .Q(n4036), .QN(n126)
         );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n3030), .CK(CLK), .Q(n4054), .QN(n133)
         );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n3029), .CK(CLK), .Q(n4072), .QN(n140)
         );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n3028), .CK(CLK), .Q(n4108), .QN(n154)
         );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n3027), .CK(CLK), .Q(n4126), .QN(n161)
         );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n3026), .CK(CLK), .Q(n4144), .QN(n168)
         );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n3025), .CK(CLK), .Q(n4162), .QN(n175)
         );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n3024), .CK(CLK), .Q(n4180), .QN(n182)
         );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n3023), .CK(CLK), .Q(n4198), .QN(n189)
         );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n3022), .CK(CLK), .Q(n4216), .QN(n196)
         );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n3021), .CK(CLK), .Q(n4234), .QN(n203)
         );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n3020), .CK(CLK), .Q(n4252), .QN(n210)
         );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n3019), .CK(CLK), .Q(n4270), .QN(n217)
         );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n3018), .CK(CLK), .Q(n3730), .QN(n7) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n3017), .CK(CLK), .Q(n3748), .QN(n14) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n3016), .CK(CLK), .Q(n3766), .QN(n21) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n3015), .CK(CLK), .Q(n3784), .QN(n28) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n3014), .CK(CLK), .Q(n3802), .QN(n35) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n3013), .CK(CLK), .Q(n3820), .QN(n42) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n3012), .CK(CLK), .Q(n3838), .QN(n49) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n3011), .CK(CLK), .Q(n3892), .QN(n70) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n3010), .CK(CLK), .Q(n4090), .QN(n147) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n3009), .CK(CLK), .Q(n4288), .QN(n224) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n3008), .CK(CLK), .Q(n3857), .QN(n280)
         );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n3007), .CK(CLK), .Q(n3875), .QN(n287)
         );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n3006), .CK(CLK), .Q(n3911), .QN(n301)
         );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n3005), .CK(CLK), .Q(n3929), .QN(n308)
         );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n3004), .CK(CLK), .Q(n3947), .QN(n315)
         );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n3003), .CK(CLK), .Q(n3965), .QN(n322)
         );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n3002), .CK(CLK), .Q(n3983), .QN(n329)
         );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n3001), .CK(CLK), .Q(n4001), .QN(n336)
         );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n3000), .CK(CLK), .Q(n4019), .QN(n343)
         );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n2999), .CK(CLK), .Q(n4037), .QN(n350)
         );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n2998), .CK(CLK), .Q(n4055), .QN(n357)
         );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n2997), .CK(CLK), .Q(n4073), .QN(n364)
         );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n2996), .CK(CLK), .Q(n4109), .QN(n378)
         );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n2995), .CK(CLK), .Q(n4127), .QN(n385)
         );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n2994), .CK(CLK), .Q(n4145), .QN(n392)
         );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n2993), .CK(CLK), .Q(n4163), .QN(n399)
         );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n2992), .CK(CLK), .Q(n4181), .QN(n406)
         );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n2991), .CK(CLK), .Q(n4199), .QN(n413)
         );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n2990), .CK(CLK), .Q(n4217), .QN(n420)
         );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n2989), .CK(CLK), .Q(n4235), .QN(n427)
         );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n2988), .CK(CLK), .Q(n4253), .QN(n434)
         );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n2987), .CK(CLK), .Q(n4271), .QN(n441)
         );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n2986), .CK(CLK), .Q(n3731), .QN(n231) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n2985), .CK(CLK), .Q(n3749), .QN(n238) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n2984), .CK(CLK), .Q(n3767), .QN(n245) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n2983), .CK(CLK), .Q(n3785), .QN(n252) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n2982), .CK(CLK), .Q(n3803), .QN(n259) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n2981), .CK(CLK), .Q(n3821), .QN(n266) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n2980), .CK(CLK), .Q(n3839), .QN(n273) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n2979), .CK(CLK), .Q(n3893), .QN(n294) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n2978), .CK(CLK), .Q(n4091), .QN(n371) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n2977), .CK(CLK), .Q(n4289), .QN(n448) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n2976), .CK(CLK), .Q(n1225) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n2975), .CK(CLK), .Q(n1227) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n2974), .CK(CLK), .Q(n1228) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n2973), .CK(CLK), .Q(n1229) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n2972), .CK(CLK), .Q(n1230) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n2971), .CK(CLK), .Q(n1231) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n2970), .CK(CLK), .Q(n1232) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n2969), .CK(CLK), .Q(n1233) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n2968), .CK(CLK), .Q(n1234) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n2967), .CK(CLK), .Q(n1235) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n2966), .CK(CLK), .Q(n1236) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n2965), .CK(CLK), .Q(n1237) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n2964), .CK(CLK), .Q(n1238) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n2963), .CK(CLK), .Q(n1239) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n2962), .CK(CLK), .Q(n1240) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n2961), .CK(CLK), .Q(n1241) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n2960), .CK(CLK), .Q(n1242) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n2959), .CK(CLK), .Q(n1243) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n2958), .CK(CLK), .Q(n1244) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n2957), .CK(CLK), .Q(n1245) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n2956), .CK(CLK), .Q(n1246) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n2955), .CK(CLK), .Q(n1247) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n2954), .CK(CLK), .Q(n1248) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n2953), .CK(CLK), .Q(n1249) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n2952), .CK(CLK), .Q(n1250) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n2951), .CK(CLK), .Q(n1251) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n2950), .CK(CLK), .Q(n1252) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n2949), .CK(CLK), .Q(n1253) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n2948), .CK(CLK), .Q(n1254) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n2947), .CK(CLK), .Q(n1255) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n2946), .CK(CLK), .Q(n1256) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n2945), .CK(CLK), .Q(n1257) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n2944), .CK(CLK), .Q(n1258) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n2943), .CK(CLK), .Q(n1260) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n2942), .CK(CLK), .Q(n1261) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n2941), .CK(CLK), .Q(n1262) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n2940), .CK(CLK), .Q(n1263) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n2939), .CK(CLK), .Q(n1264) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n2938), .CK(CLK), .Q(n1265) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n2937), .CK(CLK), .Q(n1266) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n2936), .CK(CLK), .Q(n1267) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n2935), .CK(CLK), .Q(n1268) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n2934), .CK(CLK), .Q(n1269) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n2933), .CK(CLK), .Q(n1270) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n2932), .CK(CLK), .Q(n1271) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n2931), .CK(CLK), .Q(n1272) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n2930), .CK(CLK), .Q(n1273) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n2929), .CK(CLK), .Q(n1274) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n2928), .CK(CLK), .Q(n1275) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n2927), .CK(CLK), .Q(n1276) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n2926), .CK(CLK), .Q(n1277) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n2925), .CK(CLK), .Q(n1278) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n2924), .CK(CLK), .Q(n1279) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n2923), .CK(CLK), .Q(n1280) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n2922), .CK(CLK), .Q(n1281) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n2921), .CK(CLK), .Q(n1282) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n2920), .CK(CLK), .Q(n1283) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n2919), .CK(CLK), .Q(n1284) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n2918), .CK(CLK), .Q(n1285) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n2917), .CK(CLK), .Q(n1286) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n2916), .CK(CLK), .Q(n1287) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n2915), .CK(CLK), .Q(n1288) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n2914), .CK(CLK), .Q(n1289) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n2913), .CK(CLK), .Q(n1290) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n2912), .CK(CLK), .Q(n3861), .QN(n278)
         );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n2911), .CK(CLK), .Q(n3879), .QN(n285)
         );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n2910), .CK(CLK), .Q(n3915), .QN(n299)
         );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n2909), .CK(CLK), .Q(n3933), .QN(n306)
         );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n2908), .CK(CLK), .Q(n3951), .QN(n313)
         );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n2907), .CK(CLK), .Q(n3969), .QN(n320)
         );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n2906), .CK(CLK), .Q(n3987), .QN(n327)
         );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n2905), .CK(CLK), .Q(n4005), .QN(n334)
         );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n2904), .CK(CLK), .Q(n4023), .QN(n341)
         );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n2903), .CK(CLK), .Q(n4041), .QN(n348)
         );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n2902), .CK(CLK), .Q(n4059), .QN(n355)
         );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n2901), .CK(CLK), .Q(n4077), .QN(n362)
         );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n2900), .CK(CLK), .Q(n4113), .QN(n376)
         );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n2899), .CK(CLK), .Q(n4131), .QN(n383)
         );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n2898), .CK(CLK), .Q(n4149), .QN(n390)
         );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n2897), .CK(CLK), .Q(n4167), .QN(n397)
         );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n2896), .CK(CLK), .Q(n4185), .QN(n404)
         );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n2895), .CK(CLK), .Q(n4203), .QN(n411)
         );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n2894), .CK(CLK), .Q(n4221), .QN(n418)
         );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n2893), .CK(CLK), .Q(n4239), .QN(n425)
         );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n2892), .CK(CLK), .Q(n4257), .QN(n432)
         );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n2891), .CK(CLK), .Q(n4275), .QN(n439)
         );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n2890), .CK(CLK), .Q(n3735), .QN(n229) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n2889), .CK(CLK), .Q(n3753), .QN(n236) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n2888), .CK(CLK), .Q(n3771), .QN(n243) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n2887), .CK(CLK), .Q(n3789), .QN(n250) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n2886), .CK(CLK), .Q(n3807), .QN(n257) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n2885), .CK(CLK), .Q(n3825), .QN(n264) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n2884), .CK(CLK), .Q(n3843), .QN(n271) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n2883), .CK(CLK), .Q(n3897), .QN(n292) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n2882), .CK(CLK), .Q(n4095), .QN(n369) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n2881), .CK(CLK), .Q(n4293), .QN(n446) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n2880), .CK(CLK), .Q(n3860), .QN(n54) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n2879), .CK(CLK), .Q(n3878), .QN(n61) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n2878), .CK(CLK), .Q(n3914), .QN(n75) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n2877), .CK(CLK), .Q(n3932), .QN(n82) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n2876), .CK(CLK), .Q(n3950), .QN(n89) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n2875), .CK(CLK), .Q(n3968), .QN(n96) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n2874), .CK(CLK), .Q(n3986), .QN(n103)
         );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n2873), .CK(CLK), .Q(n4004), .QN(n110)
         );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n2872), .CK(CLK), .Q(n4022), .QN(n117)
         );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n2871), .CK(CLK), .Q(n4040), .QN(n124)
         );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n2870), .CK(CLK), .Q(n4058), .QN(n131)
         );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n2869), .CK(CLK), .Q(n4076), .QN(n138)
         );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n2868), .CK(CLK), .Q(n4112), .QN(n152)
         );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n2867), .CK(CLK), .Q(n4130), .QN(n159)
         );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n2866), .CK(CLK), .Q(n4148), .QN(n166)
         );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n2865), .CK(CLK), .Q(n4166), .QN(n173)
         );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n2864), .CK(CLK), .Q(n4184), .QN(n180)
         );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n2863), .CK(CLK), .Q(n4202), .QN(n187)
         );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n2862), .CK(CLK), .Q(n4220), .QN(n194)
         );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n2861), .CK(CLK), .Q(n4238), .QN(n201)
         );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n2860), .CK(CLK), .Q(n4256), .QN(n208)
         );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n2859), .CK(CLK), .Q(n4274), .QN(n215)
         );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n2858), .CK(CLK), .Q(n3734), .QN(n5) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n2857), .CK(CLK), .Q(n3752), .QN(n12) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n2856), .CK(CLK), .Q(n3770), .QN(n19) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n2855), .CK(CLK), .Q(n3788), .QN(n26) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n2854), .CK(CLK), .Q(n3806), .QN(n33) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n2853), .CK(CLK), .Q(n3824), .QN(n40) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n2852), .CK(CLK), .Q(n3842), .QN(n47) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n2851), .CK(CLK), .Q(n3896), .QN(n68) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n2850), .CK(CLK), .Q(n4094), .QN(n145) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n2849), .CK(CLK), .Q(n4292), .QN(n222) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n2848), .CK(CLK), .Q(n1294) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n2847), .CK(CLK), .Q(n1296) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n2846), .CK(CLK), .Q(n1297) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n2845), .CK(CLK), .Q(n1298) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n2844), .CK(CLK), .Q(n1299) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n2843), .CK(CLK), .Q(n1300) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n2842), .CK(CLK), .Q(n1301) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n2841), .CK(CLK), .Q(n1302) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n2840), .CK(CLK), .Q(n1303) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n2839), .CK(CLK), .Q(n1304) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n2838), .CK(CLK), .Q(n1305) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n2837), .CK(CLK), .Q(n1306) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n2836), .CK(CLK), .Q(n1307) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n2835), .CK(CLK), .Q(n1308) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n2834), .CK(CLK), .Q(n1309) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n2833), .CK(CLK), .Q(n1310) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n2832), .CK(CLK), .Q(n1311) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n2831), .CK(CLK), .Q(n1312) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n2830), .CK(CLK), .Q(n1313) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n2829), .CK(CLK), .Q(n1314) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n2828), .CK(CLK), .Q(n1315) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2827), .CK(CLK), .Q(n1316) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n2826), .CK(CLK), .Q(n1317) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n2825), .CK(CLK), .Q(n1318) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n2824), .CK(CLK), .Q(n1319) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2823), .CK(CLK), .Q(n1320) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2822), .CK(CLK), .Q(n1321) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n2821), .CK(CLK), .Q(n1322) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2820), .CK(CLK), .Q(n1323) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n2819), .CK(CLK), .Q(n1324) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n2818), .CK(CLK), .Q(n1325) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n2817), .CK(CLK), .Q(n1326) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n2816), .CK(CLK), .Q(n1327) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n2815), .CK(CLK), .Q(n1329) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2814), .CK(CLK), .Q(n1330) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2813), .CK(CLK), .Q(n1331) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n2812), .CK(CLK), .Q(n1332) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2811), .CK(CLK), .Q(n1333) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n2810), .CK(CLK), .Q(n1334) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2809), .CK(CLK), .Q(n1335) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n2808), .CK(CLK), .Q(n1336) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2807), .CK(CLK), .Q(n1337) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n2806), .CK(CLK), .Q(n1338) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2805), .CK(CLK), .Q(n1339) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n2804), .CK(CLK), .Q(n1340) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n2803), .CK(CLK), .Q(n1341) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n2802), .CK(CLK), .Q(n1342) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n2801), .CK(CLK), .Q(n1343) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n2800), .CK(CLK), .Q(n1344) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n2799), .CK(CLK), .Q(n1345) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n2798), .CK(CLK), .Q(n1346) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n2797), .CK(CLK), .Q(n1347) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n2796), .CK(CLK), .Q(n1348) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2795), .CK(CLK), .Q(n1349) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n2794), .CK(CLK), .Q(n1350) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n2793), .CK(CLK), .Q(n1351) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n2792), .CK(CLK), .Q(n1352) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2791), .CK(CLK), .Q(n1353) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2790), .CK(CLK), .Q(n1354) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n2789), .CK(CLK), .Q(n1355) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2788), .CK(CLK), .Q(n1356) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n2787), .CK(CLK), .Q(n1357) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n2786), .CK(CLK), .Q(n1358) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n2785), .CK(CLK), .Q(n1359) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n2784), .CK(CLK), .Q(n1360), .QN(n3862)
         );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n2783), .CK(CLK), .Q(n1362), .QN(n3880)
         );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n2782), .CK(CLK), .Q(n1363), .QN(n3916)
         );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n2781), .CK(CLK), .Q(n1364), .QN(n3934)
         );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n2780), .CK(CLK), .Q(n1365), .QN(n3952)
         );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n2779), .CK(CLK), .Q(n1366), .QN(n3970)
         );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n2778), .CK(CLK), .Q(n1367), .QN(n3988)
         );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n2777), .CK(CLK), .Q(n1368), .QN(n4006)
         );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n2776), .CK(CLK), .Q(n1369), .QN(n4024)
         );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n2775), .CK(CLK), .Q(n1370), .QN(n4042)
         );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n2774), .CK(CLK), .Q(n1371), .QN(n4060)
         );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n2773), .CK(CLK), .Q(n1372), .QN(n4078)
         );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n2772), .CK(CLK), .Q(n1373), .QN(n4114)
         );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n2771), .CK(CLK), .Q(n1374), .QN(n4132)
         );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n2770), .CK(CLK), .Q(n1375), .QN(n4150)
         );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n2769), .CK(CLK), .Q(n1376), .QN(n4168)
         );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n2768), .CK(CLK), .Q(n1377), .QN(n4186)
         );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n2767), .CK(CLK), .Q(n1378), .QN(n4204)
         );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n2766), .CK(CLK), .Q(n1379), .QN(n4222)
         );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n2765), .CK(CLK), .Q(n1380), .QN(n4240)
         );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n2764), .CK(CLK), .Q(n1381), .QN(n4258)
         );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n2763), .CK(CLK), .Q(n1382), .QN(n4276)
         );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n2762), .CK(CLK), .Q(n1383), .QN(n3736)
         );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n2761), .CK(CLK), .Q(n1384), .QN(n3754)
         );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n2760), .CK(CLK), .Q(n1385), .QN(n3772)
         );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n2759), .CK(CLK), .Q(n1386), .QN(n3790)
         );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n2758), .CK(CLK), .Q(n1387), .QN(n3808)
         );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n2757), .CK(CLK), .Q(n1388), .QN(n3826)
         );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n2756), .CK(CLK), .Q(n1389), .QN(n3844)
         );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n2755), .CK(CLK), .Q(n1390), .QN(n3898)
         );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n2754), .CK(CLK), .Q(n1391), .QN(n4096)
         );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n2753), .CK(CLK), .Q(n1392), .QN(n4294)
         );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n2752), .CK(CLK), .Q(n1396), .QN(n3863)
         );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n2751), .CK(CLK), .Q(n1398), .QN(n3881)
         );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n2750), .CK(CLK), .Q(n1399), .QN(n3917)
         );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n2749), .CK(CLK), .Q(n1400), .QN(n3935)
         );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n2748), .CK(CLK), .Q(n1401), .QN(n3953)
         );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n2747), .CK(CLK), .Q(n1402), .QN(n3971)
         );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n2746), .CK(CLK), .Q(n1403), .QN(n3989)
         );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n2745), .CK(CLK), .Q(n1404), .QN(n4007)
         );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n2744), .CK(CLK), .Q(n1405), .QN(n4025)
         );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n2743), .CK(CLK), .Q(n1406), .QN(n4043)
         );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n2742), .CK(CLK), .Q(n1407), .QN(n4061)
         );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n2741), .CK(CLK), .Q(n1408), .QN(n4079)
         );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n2740), .CK(CLK), .Q(n1409), .QN(n4115)
         );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n2739), .CK(CLK), .Q(n1410), .QN(n4133)
         );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n2738), .CK(CLK), .Q(n1411), .QN(n4151)
         );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n2737), .CK(CLK), .Q(n1412), .QN(n4169)
         );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n2736), .CK(CLK), .Q(n1413), .QN(n4187)
         );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n2735), .CK(CLK), .Q(n1414), .QN(n4205)
         );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n2734), .CK(CLK), .Q(n1415), .QN(n4223)
         );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n2733), .CK(CLK), .Q(n1416), .QN(n4241)
         );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n2732), .CK(CLK), .Q(n1417), .QN(n4259)
         );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n2731), .CK(CLK), .Q(n1418), .QN(n4277)
         );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n2730), .CK(CLK), .Q(n1419), .QN(n3737)
         );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n2729), .CK(CLK), .Q(n1420), .QN(n3755)
         );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n2728), .CK(CLK), .Q(n1421), .QN(n3773)
         );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n2727), .CK(CLK), .Q(n1422), .QN(n3791)
         );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n2726), .CK(CLK), .Q(n1423), .QN(n3809)
         );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n2725), .CK(CLK), .Q(n1424), .QN(n3827)
         );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n2724), .CK(CLK), .Q(n1425), .QN(n3845)
         );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n2723), .CK(CLK), .Q(n1426), .QN(n3899)
         );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n2722), .CK(CLK), .Q(n1427), .QN(n4097)
         );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n2721), .CK(CLK), .Q(n1428), .QN(n4295)
         );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n2720), .CK(CLK), .Q(n3865) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n2719), .CK(CLK), .Q(n3883) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2718), .CK(CLK), .Q(n3919) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2717), .CK(CLK), .Q(n3937) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n2716), .CK(CLK), .Q(n3955) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2715), .CK(CLK), .Q(n3973) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n2714), .CK(CLK), .Q(n3991) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n2713), .CK(CLK), .Q(n4009) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n2712), .CK(CLK), .Q(n4027) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2711), .CK(CLK), .Q(n4045) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n2710), .CK(CLK), .Q(n4063) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2709), .CK(CLK), .Q(n4081) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n2708), .CK(CLK), .Q(n4117) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n2707), .CK(CLK), .Q(n4135) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n2706), .CK(CLK), .Q(n4153) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n2705), .CK(CLK), .Q(n4171) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n2704), .CK(CLK), .Q(n4189) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n2703), .CK(CLK), .Q(n4207) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n2702), .CK(CLK), .Q(n4225) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n2701), .CK(CLK), .Q(n4243) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n2700), .CK(CLK), .Q(n4261) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2699), .CK(CLK), .Q(n4279) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n2698), .CK(CLK), .Q(n3739) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n2697), .CK(CLK), .Q(n3757) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n2696), .CK(CLK), .Q(n3775) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2695), .CK(CLK), .Q(n3793) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2694), .CK(CLK), .Q(n3811) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n2693), .CK(CLK), .Q(n3829) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2692), .CK(CLK), .Q(n3847) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n2691), .CK(CLK), .Q(n3901) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n2690), .CK(CLK), .Q(n4099) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n2689), .CK(CLK), .Q(n4297) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n2688), .CK(CLK), .Q(n3864) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n2687), .CK(CLK), .Q(n3882) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2686), .CK(CLK), .Q(n3918) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n2685), .CK(CLK), .Q(n3936) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n2684), .CK(CLK), .Q(n3954) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2683), .CK(CLK), .Q(n3972) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n2682), .CK(CLK), .Q(n3990) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2681), .CK(CLK), .Q(n4008) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n2680), .CK(CLK), .Q(n4026) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2679), .CK(CLK), .Q(n4044) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n2678), .CK(CLK), .Q(n4062) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2677), .CK(CLK), .Q(n4080) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n2676), .CK(CLK), .Q(n4116) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n2675), .CK(CLK), .Q(n4134) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n2674), .CK(CLK), .Q(n4152) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n2673), .CK(CLK), .Q(n4170) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n2672), .CK(CLK), .Q(n4188) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n2671), .CK(CLK), .Q(n4206) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n2670), .CK(CLK), .Q(n4224) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n2669), .CK(CLK), .Q(n4242) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n2668), .CK(CLK), .Q(n4260) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2667), .CK(CLK), .Q(n4278) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n2666), .CK(CLK), .Q(n3738) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n2665), .CK(CLK), .Q(n3756) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n2664), .CK(CLK), .Q(n3774) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2663), .CK(CLK), .Q(n3792) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2662), .CK(CLK), .Q(n3810) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n2661), .CK(CLK), .Q(n3828) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2660), .CK(CLK), .Q(n3846) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n2659), .CK(CLK), .Q(n3900) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n2658), .CK(CLK), .Q(n4098) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n2657), .CK(CLK), .Q(n4296) );
  NOR3_X2 U3 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n2054), .ZN(n2031) );
  NOR3_X2 U4 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n3705), .ZN(n3682) );
  NOR3_X2 U5 ( .A1(n2056), .A2(ADD_RD2[1]), .A3(n2054), .ZN(n2034) );
  NOR3_X2 U6 ( .A1(n3707), .A2(ADD_RD1[1]), .A3(n3705), .ZN(n3685) );
  INV_X1 U7 ( .A(n835), .ZN(n833) );
  INV_X1 U8 ( .A(n835), .ZN(n834) );
  BUF_X1 U9 ( .A(n1430), .Z(n638) );
  BUF_X1 U10 ( .A(n1430), .Z(n639) );
  BUF_X1 U11 ( .A(n1429), .Z(n635) );
  BUF_X1 U12 ( .A(n1429), .Z(n636) );
  BUF_X1 U13 ( .A(n1397), .Z(n632) );
  BUF_X1 U14 ( .A(n1397), .Z(n633) );
  BUF_X1 U15 ( .A(n1361), .Z(n629) );
  BUF_X1 U16 ( .A(n1361), .Z(n630) );
  BUF_X1 U17 ( .A(n1328), .Z(n626) );
  BUF_X1 U18 ( .A(n1328), .Z(n627) );
  BUF_X1 U19 ( .A(n1295), .Z(n623) );
  BUF_X1 U20 ( .A(n1295), .Z(n624) );
  BUF_X1 U21 ( .A(n1293), .Z(n620) );
  BUF_X1 U22 ( .A(n1293), .Z(n621) );
  BUF_X1 U23 ( .A(n1291), .Z(n617) );
  BUF_X1 U24 ( .A(n1291), .Z(n618) );
  BUF_X1 U25 ( .A(n1259), .Z(n614) );
  BUF_X1 U26 ( .A(n1259), .Z(n615) );
  BUF_X1 U27 ( .A(n1226), .Z(n611) );
  BUF_X1 U28 ( .A(n1226), .Z(n612) );
  BUF_X1 U29 ( .A(n1224), .Z(n608) );
  BUF_X1 U30 ( .A(n1224), .Z(n609) );
  BUF_X1 U31 ( .A(n1222), .Z(n605) );
  BUF_X1 U32 ( .A(n1222), .Z(n606) );
  BUF_X1 U33 ( .A(n1189), .Z(n602) );
  BUF_X1 U34 ( .A(n1189), .Z(n603) );
  BUF_X1 U35 ( .A(n1156), .Z(n599) );
  BUF_X1 U36 ( .A(n1156), .Z(n600) );
  BUF_X1 U37 ( .A(n1154), .Z(n596) );
  BUF_X1 U38 ( .A(n1154), .Z(n597) );
  BUF_X1 U39 ( .A(n1152), .Z(n593) );
  BUF_X1 U40 ( .A(n1152), .Z(n594) );
  BUF_X1 U41 ( .A(n1119), .Z(n590) );
  BUF_X1 U42 ( .A(n1119), .Z(n591) );
  BUF_X1 U43 ( .A(n1086), .Z(n587) );
  BUF_X1 U44 ( .A(n1086), .Z(n588) );
  BUF_X1 U45 ( .A(n1084), .Z(n584) );
  BUF_X1 U46 ( .A(n1084), .Z(n585) );
  BUF_X1 U47 ( .A(n1082), .Z(n581) );
  BUF_X1 U48 ( .A(n1082), .Z(n582) );
  BUF_X1 U49 ( .A(n1050), .Z(n578) );
  BUF_X1 U50 ( .A(n1050), .Z(n579) );
  BUF_X1 U51 ( .A(n1017), .Z(n575) );
  BUF_X1 U52 ( .A(n1017), .Z(n576) );
  BUF_X1 U53 ( .A(n1015), .Z(n572) );
  BUF_X1 U54 ( .A(n1015), .Z(n573) );
  BUF_X1 U55 ( .A(n1013), .Z(n569) );
  BUF_X1 U56 ( .A(n1013), .Z(n570) );
  BUF_X1 U57 ( .A(n981), .Z(n566) );
  BUF_X1 U58 ( .A(n981), .Z(n567) );
  BUF_X1 U59 ( .A(n948), .Z(n563) );
  BUF_X1 U60 ( .A(n948), .Z(n564) );
  BUF_X1 U61 ( .A(n946), .Z(n560) );
  BUF_X1 U62 ( .A(n946), .Z(n561) );
  BUF_X1 U63 ( .A(n944), .Z(n557) );
  BUF_X1 U64 ( .A(n944), .Z(n558) );
  BUF_X1 U65 ( .A(n908), .Z(n554) );
  BUF_X1 U66 ( .A(n908), .Z(n555) );
  BUF_X1 U67 ( .A(n874), .Z(n551) );
  BUF_X1 U68 ( .A(n874), .Z(n552) );
  BUF_X1 U69 ( .A(n871), .Z(n548) );
  BUF_X1 U70 ( .A(n871), .Z(n549) );
  BUF_X1 U71 ( .A(n837), .Z(n452) );
  BUF_X1 U72 ( .A(n837), .Z(n453) );
  BUF_X1 U73 ( .A(n2090), .Z(n791) );
  BUF_X1 U74 ( .A(n2090), .Z(n792) );
  BUF_X1 U75 ( .A(n1464), .Z(n695) );
  BUF_X1 U76 ( .A(n1464), .Z(n696) );
  BUF_X1 U77 ( .A(n1430), .Z(n640) );
  BUF_X1 U78 ( .A(n1429), .Z(n637) );
  BUF_X1 U79 ( .A(n1397), .Z(n634) );
  BUF_X1 U80 ( .A(n1295), .Z(n625) );
  BUF_X1 U81 ( .A(n1293), .Z(n622) );
  BUF_X1 U82 ( .A(n1361), .Z(n631) );
  BUF_X1 U83 ( .A(n1328), .Z(n628) );
  BUF_X1 U84 ( .A(n1291), .Z(n619) );
  BUF_X1 U85 ( .A(n1259), .Z(n616) );
  BUF_X1 U86 ( .A(n1226), .Z(n613) );
  BUF_X1 U87 ( .A(n1224), .Z(n610) );
  BUF_X1 U88 ( .A(n1222), .Z(n607) );
  BUF_X1 U89 ( .A(n1189), .Z(n604) );
  BUF_X1 U90 ( .A(n1156), .Z(n601) );
  BUF_X1 U91 ( .A(n1154), .Z(n598) );
  BUF_X1 U92 ( .A(n1152), .Z(n595) );
  BUF_X1 U93 ( .A(n1119), .Z(n592) );
  BUF_X1 U94 ( .A(n1086), .Z(n589) );
  BUF_X1 U95 ( .A(n1084), .Z(n586) );
  BUF_X1 U96 ( .A(n1082), .Z(n583) );
  BUF_X1 U97 ( .A(n1050), .Z(n580) );
  BUF_X1 U98 ( .A(n1017), .Z(n577) );
  BUF_X1 U99 ( .A(n1015), .Z(n574) );
  BUF_X1 U100 ( .A(n946), .Z(n562) );
  BUF_X1 U101 ( .A(n1013), .Z(n571) );
  BUF_X1 U102 ( .A(n981), .Z(n568) );
  BUF_X1 U103 ( .A(n948), .Z(n565) );
  BUF_X1 U104 ( .A(n944), .Z(n559) );
  BUF_X1 U105 ( .A(n908), .Z(n556) );
  BUF_X1 U106 ( .A(n874), .Z(n553) );
  BUF_X1 U107 ( .A(n871), .Z(n550) );
  BUF_X1 U108 ( .A(n837), .Z(n454) );
  BUF_X1 U109 ( .A(n2090), .Z(n793) );
  BUF_X1 U110 ( .A(n1464), .Z(n697) );
  BUF_X1 U111 ( .A(n2076), .Z(n767) );
  BUF_X1 U112 ( .A(n2076), .Z(n768) );
  BUF_X1 U113 ( .A(n1450), .Z(n671) );
  BUF_X1 U114 ( .A(n1450), .Z(n672) );
  BUF_X1 U115 ( .A(n2095), .Z(n803) );
  BUF_X1 U116 ( .A(n2100), .Z(n815) );
  BUF_X1 U117 ( .A(n2105), .Z(n827) );
  BUF_X1 U118 ( .A(n2066), .Z(n743) );
  BUF_X1 U119 ( .A(n2071), .Z(n755) );
  BUF_X1 U120 ( .A(n2081), .Z(n779) );
  BUF_X1 U121 ( .A(n2095), .Z(n804) );
  BUF_X1 U122 ( .A(n2100), .Z(n816) );
  BUF_X1 U123 ( .A(n2105), .Z(n828) );
  BUF_X1 U124 ( .A(n2066), .Z(n744) );
  BUF_X1 U125 ( .A(n2071), .Z(n756) );
  BUF_X1 U126 ( .A(n2081), .Z(n780) );
  BUF_X1 U127 ( .A(n1455), .Z(n683) );
  BUF_X1 U128 ( .A(n1445), .Z(n659) );
  BUF_X1 U129 ( .A(n1440), .Z(n647) );
  BUF_X1 U130 ( .A(n1479), .Z(n731) );
  BUF_X1 U131 ( .A(n1469), .Z(n707) );
  BUF_X1 U132 ( .A(n1474), .Z(n719) );
  BUF_X1 U133 ( .A(n1455), .Z(n684) );
  BUF_X1 U134 ( .A(n1445), .Z(n660) );
  BUF_X1 U135 ( .A(n1440), .Z(n648) );
  BUF_X1 U136 ( .A(n1479), .Z(n732) );
  BUF_X1 U137 ( .A(n1469), .Z(n708) );
  BUF_X1 U138 ( .A(n1474), .Z(n720) );
  BUF_X1 U139 ( .A(n1442), .Z(n653) );
  BUF_X1 U140 ( .A(n1437), .Z(n641) );
  BUF_X1 U141 ( .A(n1461), .Z(n689) );
  BUF_X1 U142 ( .A(n1476), .Z(n725) );
  BUF_X1 U143 ( .A(n1466), .Z(n701) );
  BUF_X1 U144 ( .A(n1471), .Z(n713) );
  BUF_X1 U145 ( .A(n1442), .Z(n654) );
  BUF_X1 U146 ( .A(n1437), .Z(n642) );
  BUF_X1 U147 ( .A(n1461), .Z(n690) );
  BUF_X1 U148 ( .A(n1476), .Z(n726) );
  BUF_X1 U149 ( .A(n1466), .Z(n702) );
  BUF_X1 U150 ( .A(n1471), .Z(n714) );
  BUF_X1 U151 ( .A(n2087), .Z(n785) );
  BUF_X1 U152 ( .A(n2092), .Z(n797) );
  BUF_X1 U153 ( .A(n2097), .Z(n809) );
  BUF_X1 U154 ( .A(n2102), .Z(n821) );
  BUF_X1 U155 ( .A(n2063), .Z(n737) );
  BUF_X1 U156 ( .A(n2068), .Z(n749) );
  BUF_X1 U157 ( .A(n2087), .Z(n786) );
  BUF_X1 U158 ( .A(n2092), .Z(n798) );
  BUF_X1 U159 ( .A(n2097), .Z(n810) );
  BUF_X1 U160 ( .A(n2102), .Z(n822) );
  BUF_X1 U161 ( .A(n2063), .Z(n738) );
  BUF_X1 U162 ( .A(n2068), .Z(n750) );
  BUF_X1 U163 ( .A(n1452), .Z(n677) );
  BUF_X1 U164 ( .A(n1447), .Z(n665) );
  BUF_X1 U165 ( .A(n1452), .Z(n678) );
  BUF_X1 U166 ( .A(n1447), .Z(n666) );
  BUF_X1 U167 ( .A(n2073), .Z(n761) );
  BUF_X1 U168 ( .A(n2078), .Z(n773) );
  BUF_X1 U169 ( .A(n2073), .Z(n762) );
  BUF_X1 U170 ( .A(n2078), .Z(n774) );
  BUF_X1 U171 ( .A(n1443), .Z(n656) );
  BUF_X1 U172 ( .A(n1438), .Z(n644) );
  BUF_X1 U173 ( .A(n1462), .Z(n692) );
  BUF_X1 U174 ( .A(n1477), .Z(n728) );
  BUF_X1 U175 ( .A(n1467), .Z(n704) );
  BUF_X1 U176 ( .A(n1472), .Z(n716) );
  BUF_X1 U177 ( .A(n1443), .Z(n657) );
  BUF_X1 U178 ( .A(n1438), .Z(n645) );
  BUF_X1 U179 ( .A(n1462), .Z(n693) );
  BUF_X1 U180 ( .A(n1477), .Z(n729) );
  BUF_X1 U181 ( .A(n1467), .Z(n705) );
  BUF_X1 U182 ( .A(n1472), .Z(n717) );
  BUF_X1 U183 ( .A(n2088), .Z(n788) );
  BUF_X1 U184 ( .A(n2093), .Z(n800) );
  BUF_X1 U185 ( .A(n2098), .Z(n812) );
  BUF_X1 U186 ( .A(n2103), .Z(n824) );
  BUF_X1 U187 ( .A(n2064), .Z(n740) );
  BUF_X1 U188 ( .A(n2069), .Z(n752) );
  BUF_X1 U189 ( .A(n2088), .Z(n789) );
  BUF_X1 U190 ( .A(n2093), .Z(n801) );
  BUF_X1 U191 ( .A(n2098), .Z(n813) );
  BUF_X1 U192 ( .A(n2103), .Z(n825) );
  BUF_X1 U193 ( .A(n2064), .Z(n741) );
  BUF_X1 U194 ( .A(n2069), .Z(n753) );
  BUF_X1 U195 ( .A(n2077), .Z(n770) );
  BUF_X1 U196 ( .A(n2077), .Z(n771) );
  BUF_X1 U197 ( .A(n1451), .Z(n674) );
  BUF_X1 U198 ( .A(n1451), .Z(n675) );
  BUF_X1 U199 ( .A(n1453), .Z(n680) );
  BUF_X1 U200 ( .A(n1448), .Z(n668) );
  BUF_X1 U201 ( .A(n1453), .Z(n681) );
  BUF_X1 U202 ( .A(n1448), .Z(n669) );
  BUF_X1 U203 ( .A(n2091), .Z(n794) );
  BUF_X1 U204 ( .A(n2096), .Z(n806) );
  BUF_X1 U205 ( .A(n2101), .Z(n818) );
  BUF_X1 U206 ( .A(n2106), .Z(n830) );
  BUF_X1 U207 ( .A(n2067), .Z(n746) );
  BUF_X1 U208 ( .A(n2072), .Z(n758) );
  BUF_X1 U209 ( .A(n2082), .Z(n782) );
  BUF_X1 U210 ( .A(n2091), .Z(n795) );
  BUF_X1 U211 ( .A(n2096), .Z(n807) );
  BUF_X1 U212 ( .A(n2101), .Z(n819) );
  BUF_X1 U213 ( .A(n2106), .Z(n831) );
  BUF_X1 U214 ( .A(n2067), .Z(n747) );
  BUF_X1 U215 ( .A(n2072), .Z(n759) );
  BUF_X1 U216 ( .A(n2082), .Z(n783) );
  BUF_X1 U217 ( .A(n1456), .Z(n686) );
  BUF_X1 U218 ( .A(n1446), .Z(n662) );
  BUF_X1 U219 ( .A(n1441), .Z(n650) );
  BUF_X1 U220 ( .A(n1465), .Z(n698) );
  BUF_X1 U221 ( .A(n1480), .Z(n734) );
  BUF_X1 U222 ( .A(n1470), .Z(n710) );
  BUF_X1 U223 ( .A(n1475), .Z(n722) );
  BUF_X1 U224 ( .A(n1456), .Z(n687) );
  BUF_X1 U225 ( .A(n1446), .Z(n663) );
  BUF_X1 U226 ( .A(n1441), .Z(n651) );
  BUF_X1 U227 ( .A(n1465), .Z(n699) );
  BUF_X1 U228 ( .A(n1480), .Z(n735) );
  BUF_X1 U229 ( .A(n1470), .Z(n711) );
  BUF_X1 U230 ( .A(n1475), .Z(n723) );
  BUF_X1 U231 ( .A(n2074), .Z(n764) );
  BUF_X1 U232 ( .A(n2079), .Z(n776) );
  BUF_X1 U233 ( .A(n2074), .Z(n765) );
  BUF_X1 U234 ( .A(n2079), .Z(n777) );
  BUF_X1 U235 ( .A(n2076), .Z(n769) );
  BUF_X1 U236 ( .A(n1450), .Z(n673) );
  BUF_X1 U237 ( .A(n2095), .Z(n805) );
  BUF_X1 U238 ( .A(n2100), .Z(n817) );
  BUF_X1 U239 ( .A(n2105), .Z(n829) );
  BUF_X1 U240 ( .A(n2066), .Z(n745) );
  BUF_X1 U241 ( .A(n2071), .Z(n757) );
  BUF_X1 U242 ( .A(n2081), .Z(n781) );
  BUF_X1 U243 ( .A(n1455), .Z(n685) );
  BUF_X1 U244 ( .A(n1445), .Z(n661) );
  BUF_X1 U245 ( .A(n1440), .Z(n649) );
  BUF_X1 U246 ( .A(n1479), .Z(n733) );
  BUF_X1 U247 ( .A(n1469), .Z(n709) );
  BUF_X1 U248 ( .A(n1474), .Z(n721) );
  BUF_X1 U249 ( .A(n1442), .Z(n655) );
  BUF_X1 U250 ( .A(n1437), .Z(n643) );
  BUF_X1 U251 ( .A(n1461), .Z(n691) );
  BUF_X1 U252 ( .A(n1476), .Z(n727) );
  BUF_X1 U253 ( .A(n1466), .Z(n703) );
  BUF_X1 U254 ( .A(n1471), .Z(n715) );
  BUF_X1 U255 ( .A(n2087), .Z(n787) );
  BUF_X1 U256 ( .A(n2092), .Z(n799) );
  BUF_X1 U257 ( .A(n2097), .Z(n811) );
  BUF_X1 U258 ( .A(n2102), .Z(n823) );
  BUF_X1 U259 ( .A(n2063), .Z(n739) );
  BUF_X1 U260 ( .A(n2068), .Z(n751) );
  BUF_X1 U261 ( .A(n1452), .Z(n679) );
  BUF_X1 U262 ( .A(n1447), .Z(n667) );
  BUF_X1 U263 ( .A(n2073), .Z(n763) );
  BUF_X1 U264 ( .A(n2078), .Z(n775) );
  BUF_X1 U265 ( .A(n1443), .Z(n658) );
  BUF_X1 U266 ( .A(n1438), .Z(n646) );
  BUF_X1 U267 ( .A(n1462), .Z(n694) );
  BUF_X1 U268 ( .A(n1477), .Z(n730) );
  BUF_X1 U269 ( .A(n1467), .Z(n706) );
  BUF_X1 U270 ( .A(n1472), .Z(n718) );
  BUF_X1 U271 ( .A(n2088), .Z(n790) );
  BUF_X1 U272 ( .A(n2093), .Z(n802) );
  BUF_X1 U273 ( .A(n2098), .Z(n814) );
  BUF_X1 U274 ( .A(n2103), .Z(n826) );
  BUF_X1 U275 ( .A(n2064), .Z(n742) );
  BUF_X1 U276 ( .A(n2069), .Z(n754) );
  BUF_X1 U277 ( .A(n2077), .Z(n772) );
  BUF_X1 U278 ( .A(n1451), .Z(n676) );
  BUF_X1 U279 ( .A(n1453), .Z(n682) );
  BUF_X1 U280 ( .A(n1448), .Z(n670) );
  BUF_X1 U281 ( .A(n2074), .Z(n766) );
  BUF_X1 U282 ( .A(n2079), .Z(n778) );
  BUF_X1 U283 ( .A(n2091), .Z(n796) );
  BUF_X1 U284 ( .A(n2106), .Z(n832) );
  BUF_X1 U285 ( .A(n2072), .Z(n760) );
  BUF_X1 U286 ( .A(n2082), .Z(n784) );
  BUF_X1 U287 ( .A(n1456), .Z(n688) );
  BUF_X1 U288 ( .A(n1446), .Z(n664) );
  BUF_X1 U289 ( .A(n1465), .Z(n700) );
  BUF_X1 U290 ( .A(n1480), .Z(n736) );
  BUF_X1 U291 ( .A(n2096), .Z(n808) );
  BUF_X1 U292 ( .A(n2101), .Z(n820) );
  BUF_X1 U293 ( .A(n2067), .Z(n748) );
  BUF_X1 U294 ( .A(n1441), .Z(n652) );
  BUF_X1 U295 ( .A(n1470), .Z(n712) );
  BUF_X1 U296 ( .A(n1475), .Z(n724) );
  BUF_X1 U297 ( .A(n868), .Z(n546) );
  BUF_X1 U298 ( .A(n867), .Z(n543) );
  BUF_X1 U299 ( .A(n866), .Z(n540) );
  BUF_X1 U300 ( .A(n865), .Z(n537) );
  BUF_X1 U301 ( .A(n864), .Z(n534) );
  BUF_X1 U302 ( .A(n863), .Z(n531) );
  BUF_X1 U303 ( .A(n862), .Z(n528) );
  BUF_X1 U304 ( .A(n861), .Z(n525) );
  BUF_X1 U305 ( .A(n860), .Z(n522) );
  BUF_X1 U306 ( .A(n859), .Z(n519) );
  BUF_X1 U307 ( .A(n858), .Z(n516) );
  BUF_X1 U308 ( .A(n857), .Z(n513) );
  BUF_X1 U309 ( .A(n856), .Z(n510) );
  BUF_X1 U310 ( .A(n855), .Z(n507) );
  BUF_X1 U311 ( .A(n854), .Z(n504) );
  BUF_X1 U312 ( .A(n853), .Z(n501) );
  BUF_X1 U313 ( .A(n852), .Z(n498) );
  BUF_X1 U314 ( .A(n851), .Z(n495) );
  BUF_X1 U315 ( .A(n850), .Z(n492) );
  BUF_X1 U316 ( .A(n849), .Z(n489) );
  BUF_X1 U317 ( .A(n848), .Z(n486) );
  BUF_X1 U318 ( .A(n847), .Z(n483) );
  BUF_X1 U319 ( .A(n846), .Z(n480) );
  BUF_X1 U320 ( .A(n845), .Z(n477) );
  BUF_X1 U321 ( .A(n844), .Z(n474) );
  BUF_X1 U322 ( .A(n843), .Z(n471) );
  BUF_X1 U323 ( .A(n842), .Z(n468) );
  BUF_X1 U324 ( .A(n841), .Z(n465) );
  BUF_X1 U325 ( .A(n840), .Z(n462) );
  BUF_X1 U326 ( .A(n839), .Z(n459) );
  BUF_X1 U327 ( .A(n838), .Z(n456) );
  BUF_X1 U328 ( .A(n836), .Z(n450) );
  BUF_X1 U329 ( .A(n868), .Z(n545) );
  BUF_X1 U330 ( .A(n867), .Z(n542) );
  BUF_X1 U331 ( .A(n866), .Z(n539) );
  BUF_X1 U332 ( .A(n865), .Z(n536) );
  BUF_X1 U333 ( .A(n864), .Z(n533) );
  BUF_X1 U334 ( .A(n863), .Z(n530) );
  BUF_X1 U335 ( .A(n862), .Z(n527) );
  BUF_X1 U336 ( .A(n861), .Z(n524) );
  BUF_X1 U337 ( .A(n860), .Z(n521) );
  BUF_X1 U338 ( .A(n859), .Z(n518) );
  BUF_X1 U339 ( .A(n858), .Z(n515) );
  BUF_X1 U340 ( .A(n857), .Z(n512) );
  BUF_X1 U341 ( .A(n856), .Z(n509) );
  BUF_X1 U342 ( .A(n855), .Z(n506) );
  BUF_X1 U343 ( .A(n854), .Z(n503) );
  BUF_X1 U344 ( .A(n853), .Z(n500) );
  BUF_X1 U345 ( .A(n852), .Z(n497) );
  BUF_X1 U346 ( .A(n851), .Z(n494) );
  BUF_X1 U347 ( .A(n850), .Z(n491) );
  BUF_X1 U348 ( .A(n849), .Z(n488) );
  BUF_X1 U349 ( .A(n848), .Z(n485) );
  BUF_X1 U350 ( .A(n847), .Z(n482) );
  BUF_X1 U351 ( .A(n846), .Z(n479) );
  BUF_X1 U352 ( .A(n845), .Z(n476) );
  BUF_X1 U353 ( .A(n844), .Z(n473) );
  BUF_X1 U354 ( .A(n843), .Z(n470) );
  BUF_X1 U355 ( .A(n842), .Z(n467) );
  BUF_X1 U356 ( .A(n841), .Z(n464) );
  BUF_X1 U357 ( .A(n840), .Z(n461) );
  BUF_X1 U358 ( .A(n839), .Z(n458) );
  BUF_X1 U359 ( .A(n838), .Z(n455) );
  BUF_X1 U360 ( .A(n836), .Z(n449) );
  BUF_X1 U361 ( .A(n868), .Z(n547) );
  BUF_X1 U362 ( .A(n839), .Z(n460) );
  BUF_X1 U363 ( .A(n836), .Z(n451) );
  BUF_X1 U364 ( .A(n867), .Z(n544) );
  BUF_X1 U365 ( .A(n866), .Z(n541) );
  BUF_X1 U366 ( .A(n865), .Z(n538) );
  BUF_X1 U367 ( .A(n864), .Z(n535) );
  BUF_X1 U368 ( .A(n863), .Z(n532) );
  BUF_X1 U369 ( .A(n862), .Z(n529) );
  BUF_X1 U370 ( .A(n861), .Z(n526) );
  BUF_X1 U371 ( .A(n860), .Z(n523) );
  BUF_X1 U372 ( .A(n859), .Z(n520) );
  BUF_X1 U373 ( .A(n858), .Z(n517) );
  BUF_X1 U374 ( .A(n857), .Z(n514) );
  BUF_X1 U375 ( .A(n856), .Z(n511) );
  BUF_X1 U376 ( .A(n855), .Z(n508) );
  BUF_X1 U377 ( .A(n854), .Z(n505) );
  BUF_X1 U378 ( .A(n853), .Z(n502) );
  BUF_X1 U379 ( .A(n852), .Z(n499) );
  BUF_X1 U380 ( .A(n851), .Z(n496) );
  BUF_X1 U381 ( .A(n850), .Z(n493) );
  BUF_X1 U382 ( .A(n849), .Z(n490) );
  BUF_X1 U383 ( .A(n848), .Z(n487) );
  BUF_X1 U384 ( .A(n847), .Z(n484) );
  BUF_X1 U385 ( .A(n846), .Z(n481) );
  BUF_X1 U386 ( .A(n845), .Z(n478) );
  BUF_X1 U387 ( .A(n844), .Z(n475) );
  BUF_X1 U388 ( .A(n843), .Z(n472) );
  BUF_X1 U389 ( .A(n842), .Z(n469) );
  BUF_X1 U390 ( .A(n841), .Z(n466) );
  BUF_X1 U391 ( .A(n840), .Z(n463) );
  BUF_X1 U392 ( .A(n838), .Z(n457) );
  INV_X1 U393 ( .A(RESET), .ZN(n835) );
  MUX2_X1 U394 ( .A(n3855), .B(n449), .S(n454), .Z(n3680) );
  MUX2_X1 U395 ( .A(n3873), .B(n455), .S(n454), .Z(n3679) );
  MUX2_X1 U396 ( .A(n3909), .B(n458), .S(n454), .Z(n3678) );
  MUX2_X1 U397 ( .A(n3927), .B(n461), .S(n454), .Z(n3677) );
  MUX2_X1 U398 ( .A(n3945), .B(n464), .S(n454), .Z(n3676) );
  MUX2_X1 U399 ( .A(n3963), .B(n467), .S(n454), .Z(n3675) );
  MUX2_X1 U400 ( .A(n3981), .B(n470), .S(n454), .Z(n3674) );
  MUX2_X1 U401 ( .A(n3999), .B(n473), .S(n454), .Z(n3673) );
  MUX2_X1 U402 ( .A(n4017), .B(n476), .S(n453), .Z(n3672) );
  MUX2_X1 U403 ( .A(n4035), .B(n479), .S(n453), .Z(n3671) );
  MUX2_X1 U404 ( .A(n4053), .B(n482), .S(n453), .Z(n3670) );
  MUX2_X1 U405 ( .A(n4071), .B(n485), .S(n453), .Z(n3669) );
  MUX2_X1 U406 ( .A(n4107), .B(n488), .S(n453), .Z(n3668) );
  MUX2_X1 U407 ( .A(n4125), .B(n491), .S(n453), .Z(n3667) );
  MUX2_X1 U408 ( .A(n4143), .B(n494), .S(n453), .Z(n3666) );
  MUX2_X1 U409 ( .A(n4161), .B(n497), .S(n453), .Z(n3665) );
  MUX2_X1 U410 ( .A(n4179), .B(n500), .S(n453), .Z(n3664) );
  MUX2_X1 U411 ( .A(n4197), .B(n503), .S(n453), .Z(n3663) );
  MUX2_X1 U412 ( .A(n4215), .B(n506), .S(n453), .Z(n3662) );
  MUX2_X1 U413 ( .A(n4233), .B(n509), .S(n453), .Z(n3661) );
  MUX2_X1 U414 ( .A(n4251), .B(n512), .S(n452), .Z(n3660) );
  MUX2_X1 U415 ( .A(n4269), .B(n515), .S(n452), .Z(n3659) );
  MUX2_X1 U416 ( .A(n3729), .B(n518), .S(n452), .Z(n3658) );
  MUX2_X1 U417 ( .A(n3747), .B(n521), .S(n452), .Z(n3657) );
  MUX2_X1 U418 ( .A(n3765), .B(n524), .S(n452), .Z(n3656) );
  MUX2_X1 U419 ( .A(n3783), .B(n527), .S(n452), .Z(n3655) );
  MUX2_X1 U420 ( .A(n3801), .B(n530), .S(n452), .Z(n3654) );
  MUX2_X1 U421 ( .A(n3819), .B(n533), .S(n452), .Z(n3653) );
  MUX2_X1 U422 ( .A(n3837), .B(n536), .S(n452), .Z(n3652) );
  MUX2_X1 U423 ( .A(n3891), .B(n539), .S(n452), .Z(n3651) );
  MUX2_X1 U424 ( .A(n4089), .B(n542), .S(n452), .Z(n3650) );
  MUX2_X1 U425 ( .A(n4287), .B(n545), .S(n452), .Z(n3649) );
  OAI21_X1 U426 ( .B1(n869), .B2(n870), .A(n833), .ZN(n837) );
  MUX2_X1 U427 ( .A(n3854), .B(n449), .S(n550), .Z(n3648) );
  MUX2_X1 U428 ( .A(n3872), .B(n455), .S(n550), .Z(n3647) );
  MUX2_X1 U429 ( .A(n3908), .B(n458), .S(n550), .Z(n3646) );
  MUX2_X1 U430 ( .A(n3926), .B(n461), .S(n550), .Z(n3645) );
  MUX2_X1 U431 ( .A(n3944), .B(n464), .S(n550), .Z(n3644) );
  MUX2_X1 U432 ( .A(n3962), .B(n467), .S(n550), .Z(n3643) );
  MUX2_X1 U433 ( .A(n3980), .B(n470), .S(n550), .Z(n3642) );
  MUX2_X1 U434 ( .A(n3998), .B(n473), .S(n550), .Z(n3641) );
  MUX2_X1 U435 ( .A(n4016), .B(n476), .S(n549), .Z(n3640) );
  MUX2_X1 U436 ( .A(n4034), .B(n479), .S(n549), .Z(n3639) );
  MUX2_X1 U437 ( .A(n4052), .B(n482), .S(n549), .Z(n3638) );
  MUX2_X1 U438 ( .A(n4070), .B(n485), .S(n549), .Z(n3637) );
  MUX2_X1 U439 ( .A(n4106), .B(n488), .S(n549), .Z(n3636) );
  MUX2_X1 U440 ( .A(n4124), .B(n491), .S(n549), .Z(n3635) );
  MUX2_X1 U441 ( .A(n4142), .B(n494), .S(n549), .Z(n3634) );
  MUX2_X1 U442 ( .A(n4160), .B(n497), .S(n549), .Z(n3633) );
  MUX2_X1 U443 ( .A(n4178), .B(n500), .S(n549), .Z(n3632) );
  MUX2_X1 U444 ( .A(n4196), .B(n503), .S(n549), .Z(n3631) );
  MUX2_X1 U445 ( .A(n4214), .B(n506), .S(n549), .Z(n3630) );
  MUX2_X1 U446 ( .A(n4232), .B(n509), .S(n549), .Z(n3629) );
  MUX2_X1 U447 ( .A(n4250), .B(n512), .S(n548), .Z(n3628) );
  MUX2_X1 U448 ( .A(n4268), .B(n515), .S(n548), .Z(n3627) );
  MUX2_X1 U449 ( .A(n3728), .B(n518), .S(n548), .Z(n3626) );
  MUX2_X1 U450 ( .A(n3746), .B(n521), .S(n548), .Z(n3625) );
  MUX2_X1 U451 ( .A(n3764), .B(n524), .S(n548), .Z(n3624) );
  MUX2_X1 U452 ( .A(n3782), .B(n527), .S(n548), .Z(n3623) );
  MUX2_X1 U453 ( .A(n3800), .B(n530), .S(n548), .Z(n3622) );
  MUX2_X1 U454 ( .A(n3818), .B(n533), .S(n548), .Z(n3621) );
  MUX2_X1 U455 ( .A(n3836), .B(n536), .S(n548), .Z(n3620) );
  MUX2_X1 U456 ( .A(n3890), .B(n539), .S(n548), .Z(n3619) );
  MUX2_X1 U457 ( .A(n4088), .B(n542), .S(n548), .Z(n3618) );
  MUX2_X1 U458 ( .A(n4286), .B(n545), .S(n548), .Z(n3617) );
  OAI21_X1 U459 ( .B1(n869), .B2(n872), .A(n833), .ZN(n871) );
  MUX2_X1 U460 ( .A(n873), .B(n449), .S(n553), .Z(n3616) );
  MUX2_X1 U461 ( .A(n875), .B(n455), .S(n553), .Z(n3615) );
  MUX2_X1 U462 ( .A(n876), .B(n458), .S(n553), .Z(n3614) );
  MUX2_X1 U463 ( .A(n877), .B(n461), .S(n553), .Z(n3613) );
  MUX2_X1 U464 ( .A(n878), .B(n464), .S(n553), .Z(n3612) );
  MUX2_X1 U465 ( .A(n879), .B(n467), .S(n553), .Z(n3611) );
  MUX2_X1 U466 ( .A(n880), .B(n470), .S(n553), .Z(n3610) );
  MUX2_X1 U467 ( .A(n881), .B(n473), .S(n553), .Z(n3609) );
  MUX2_X1 U468 ( .A(n882), .B(n476), .S(n552), .Z(n3608) );
  MUX2_X1 U469 ( .A(n883), .B(n479), .S(n552), .Z(n3607) );
  MUX2_X1 U470 ( .A(n884), .B(n482), .S(n552), .Z(n3606) );
  MUX2_X1 U471 ( .A(n885), .B(n485), .S(n552), .Z(n3605) );
  MUX2_X1 U472 ( .A(n886), .B(n488), .S(n552), .Z(n3604) );
  MUX2_X1 U473 ( .A(n887), .B(n491), .S(n552), .Z(n3603) );
  MUX2_X1 U474 ( .A(n888), .B(n494), .S(n552), .Z(n3602) );
  MUX2_X1 U475 ( .A(n889), .B(n497), .S(n552), .Z(n3601) );
  MUX2_X1 U476 ( .A(n890), .B(n500), .S(n552), .Z(n3600) );
  MUX2_X1 U477 ( .A(n891), .B(n503), .S(n552), .Z(n3599) );
  MUX2_X1 U478 ( .A(n892), .B(n506), .S(n552), .Z(n3598) );
  MUX2_X1 U479 ( .A(n893), .B(n509), .S(n552), .Z(n3597) );
  MUX2_X1 U480 ( .A(n894), .B(n512), .S(n551), .Z(n3596) );
  MUX2_X1 U481 ( .A(n895), .B(n515), .S(n551), .Z(n3595) );
  MUX2_X1 U482 ( .A(n896), .B(n518), .S(n551), .Z(n3594) );
  MUX2_X1 U483 ( .A(n897), .B(n521), .S(n551), .Z(n3593) );
  MUX2_X1 U484 ( .A(n898), .B(n524), .S(n551), .Z(n3592) );
  MUX2_X1 U485 ( .A(n899), .B(n527), .S(n551), .Z(n3591) );
  MUX2_X1 U486 ( .A(n900), .B(n530), .S(n551), .Z(n3590) );
  MUX2_X1 U487 ( .A(n901), .B(n533), .S(n551), .Z(n3589) );
  MUX2_X1 U488 ( .A(n902), .B(n536), .S(n551), .Z(n3588) );
  MUX2_X1 U489 ( .A(n903), .B(n539), .S(n551), .Z(n3587) );
  MUX2_X1 U490 ( .A(n904), .B(n542), .S(n551), .Z(n3586) );
  MUX2_X1 U491 ( .A(n905), .B(n545), .S(n551), .Z(n3585) );
  OAI21_X1 U492 ( .B1(n869), .B2(n906), .A(n833), .ZN(n874) );
  MUX2_X1 U493 ( .A(n907), .B(n449), .S(n556), .Z(n3584) );
  MUX2_X1 U494 ( .A(n909), .B(n455), .S(n556), .Z(n3583) );
  MUX2_X1 U495 ( .A(n910), .B(n458), .S(n556), .Z(n3582) );
  MUX2_X1 U496 ( .A(n911), .B(n461), .S(n556), .Z(n3581) );
  MUX2_X1 U497 ( .A(n912), .B(n464), .S(n556), .Z(n3580) );
  MUX2_X1 U498 ( .A(n913), .B(n467), .S(n556), .Z(n3579) );
  MUX2_X1 U499 ( .A(n914), .B(n470), .S(n556), .Z(n3578) );
  MUX2_X1 U500 ( .A(n915), .B(n473), .S(n556), .Z(n3577) );
  MUX2_X1 U501 ( .A(n916), .B(n476), .S(n555), .Z(n3576) );
  MUX2_X1 U502 ( .A(n917), .B(n479), .S(n555), .Z(n3575) );
  MUX2_X1 U503 ( .A(n918), .B(n482), .S(n555), .Z(n3574) );
  MUX2_X1 U504 ( .A(n919), .B(n485), .S(n555), .Z(n3573) );
  MUX2_X1 U505 ( .A(n920), .B(n488), .S(n555), .Z(n3572) );
  MUX2_X1 U506 ( .A(n921), .B(n491), .S(n555), .Z(n3571) );
  MUX2_X1 U507 ( .A(n922), .B(n494), .S(n555), .Z(n3570) );
  MUX2_X1 U508 ( .A(n923), .B(n497), .S(n555), .Z(n3569) );
  MUX2_X1 U509 ( .A(n924), .B(n500), .S(n555), .Z(n3568) );
  MUX2_X1 U510 ( .A(n925), .B(n503), .S(n555), .Z(n3567) );
  MUX2_X1 U511 ( .A(n926), .B(n506), .S(n555), .Z(n3566) );
  MUX2_X1 U512 ( .A(n927), .B(n509), .S(n555), .Z(n3565) );
  MUX2_X1 U513 ( .A(n928), .B(n512), .S(n554), .Z(n3564) );
  MUX2_X1 U514 ( .A(n929), .B(n515), .S(n554), .Z(n3563) );
  MUX2_X1 U515 ( .A(n930), .B(n518), .S(n554), .Z(n3562) );
  MUX2_X1 U516 ( .A(n931), .B(n521), .S(n554), .Z(n3561) );
  MUX2_X1 U517 ( .A(n932), .B(n524), .S(n554), .Z(n3560) );
  MUX2_X1 U518 ( .A(n933), .B(n527), .S(n554), .Z(n3559) );
  MUX2_X1 U519 ( .A(n934), .B(n530), .S(n554), .Z(n3558) );
  MUX2_X1 U520 ( .A(n935), .B(n533), .S(n554), .Z(n3557) );
  MUX2_X1 U521 ( .A(n936), .B(n536), .S(n554), .Z(n3556) );
  MUX2_X1 U522 ( .A(n937), .B(n539), .S(n554), .Z(n3555) );
  MUX2_X1 U523 ( .A(n938), .B(n542), .S(n554), .Z(n3554) );
  MUX2_X1 U524 ( .A(n939), .B(n545), .S(n554), .Z(n3553) );
  OAI21_X1 U525 ( .B1(n869), .B2(n940), .A(n833), .ZN(n908) );
  NAND3_X1 U526 ( .A1(n941), .A2(n942), .A3(n943), .ZN(n869) );
  MUX2_X1 U527 ( .A(n3853), .B(n449), .S(n559), .Z(n3552) );
  MUX2_X1 U528 ( .A(n3871), .B(n455), .S(n559), .Z(n3551) );
  MUX2_X1 U529 ( .A(n3907), .B(n458), .S(n559), .Z(n3550) );
  MUX2_X1 U530 ( .A(n3925), .B(n461), .S(n559), .Z(n3549) );
  MUX2_X1 U531 ( .A(n3943), .B(n464), .S(n559), .Z(n3548) );
  MUX2_X1 U532 ( .A(n3961), .B(n467), .S(n559), .Z(n3547) );
  MUX2_X1 U533 ( .A(n3979), .B(n470), .S(n559), .Z(n3546) );
  MUX2_X1 U534 ( .A(n3997), .B(n473), .S(n559), .Z(n3545) );
  MUX2_X1 U535 ( .A(n4015), .B(n476), .S(n558), .Z(n3544) );
  MUX2_X1 U536 ( .A(n4033), .B(n479), .S(n558), .Z(n3543) );
  MUX2_X1 U537 ( .A(n4051), .B(n482), .S(n558), .Z(n3542) );
  MUX2_X1 U538 ( .A(n4069), .B(n485), .S(n558), .Z(n3541) );
  MUX2_X1 U539 ( .A(n4105), .B(n488), .S(n558), .Z(n3540) );
  MUX2_X1 U540 ( .A(n4123), .B(n491), .S(n558), .Z(n3539) );
  MUX2_X1 U541 ( .A(n4141), .B(n494), .S(n558), .Z(n3538) );
  MUX2_X1 U542 ( .A(n4159), .B(n497), .S(n558), .Z(n3537) );
  MUX2_X1 U543 ( .A(n4177), .B(n500), .S(n558), .Z(n3536) );
  MUX2_X1 U544 ( .A(n4195), .B(n503), .S(n558), .Z(n3535) );
  MUX2_X1 U545 ( .A(n4213), .B(n506), .S(n558), .Z(n3534) );
  MUX2_X1 U546 ( .A(n4231), .B(n509), .S(n558), .Z(n3533) );
  MUX2_X1 U547 ( .A(n4249), .B(n512), .S(n557), .Z(n3532) );
  MUX2_X1 U548 ( .A(n4267), .B(n515), .S(n557), .Z(n3531) );
  MUX2_X1 U549 ( .A(n3727), .B(n518), .S(n557), .Z(n3530) );
  MUX2_X1 U550 ( .A(n3745), .B(n521), .S(n557), .Z(n3529) );
  MUX2_X1 U551 ( .A(n3763), .B(n524), .S(n557), .Z(n3528) );
  MUX2_X1 U552 ( .A(n3781), .B(n527), .S(n557), .Z(n3527) );
  MUX2_X1 U553 ( .A(n3799), .B(n530), .S(n557), .Z(n3526) );
  MUX2_X1 U554 ( .A(n3817), .B(n533), .S(n557), .Z(n3525) );
  MUX2_X1 U555 ( .A(n3835), .B(n536), .S(n557), .Z(n3524) );
  MUX2_X1 U556 ( .A(n3889), .B(n539), .S(n557), .Z(n3523) );
  MUX2_X1 U557 ( .A(n4087), .B(n542), .S(n557), .Z(n3522) );
  MUX2_X1 U558 ( .A(n4285), .B(n545), .S(n557), .Z(n3521) );
  OAI21_X1 U559 ( .B1(n870), .B2(n945), .A(n833), .ZN(n944) );
  MUX2_X1 U560 ( .A(n3852), .B(n449), .S(n562), .Z(n3520) );
  MUX2_X1 U561 ( .A(n3870), .B(n455), .S(n562), .Z(n3519) );
  MUX2_X1 U562 ( .A(n3906), .B(n458), .S(n562), .Z(n3518) );
  MUX2_X1 U563 ( .A(n3924), .B(n461), .S(n562), .Z(n3517) );
  MUX2_X1 U564 ( .A(n3942), .B(n464), .S(n562), .Z(n3516) );
  MUX2_X1 U565 ( .A(n3960), .B(n467), .S(n562), .Z(n3515) );
  MUX2_X1 U566 ( .A(n3978), .B(n470), .S(n562), .Z(n3514) );
  MUX2_X1 U567 ( .A(n3996), .B(n473), .S(n562), .Z(n3513) );
  MUX2_X1 U568 ( .A(n4014), .B(n476), .S(n561), .Z(n3512) );
  MUX2_X1 U569 ( .A(n4032), .B(n479), .S(n561), .Z(n3511) );
  MUX2_X1 U570 ( .A(n4050), .B(n482), .S(n561), .Z(n3510) );
  MUX2_X1 U571 ( .A(n4068), .B(n485), .S(n561), .Z(n3509) );
  MUX2_X1 U572 ( .A(n4104), .B(n488), .S(n561), .Z(n3508) );
  MUX2_X1 U573 ( .A(n4122), .B(n491), .S(n561), .Z(n3507) );
  MUX2_X1 U574 ( .A(n4140), .B(n494), .S(n561), .Z(n3506) );
  MUX2_X1 U575 ( .A(n4158), .B(n497), .S(n561), .Z(n3505) );
  MUX2_X1 U576 ( .A(n4176), .B(n500), .S(n561), .Z(n3504) );
  MUX2_X1 U577 ( .A(n4194), .B(n503), .S(n561), .Z(n3503) );
  MUX2_X1 U578 ( .A(n4212), .B(n506), .S(n561), .Z(n3502) );
  MUX2_X1 U579 ( .A(n4230), .B(n509), .S(n561), .Z(n3501) );
  MUX2_X1 U580 ( .A(n4248), .B(n512), .S(n560), .Z(n3500) );
  MUX2_X1 U581 ( .A(n4266), .B(n515), .S(n560), .Z(n3499) );
  MUX2_X1 U582 ( .A(n3726), .B(n518), .S(n560), .Z(n3498) );
  MUX2_X1 U583 ( .A(n3744), .B(n521), .S(n560), .Z(n3497) );
  MUX2_X1 U584 ( .A(n3762), .B(n524), .S(n560), .Z(n3496) );
  MUX2_X1 U585 ( .A(n3780), .B(n527), .S(n560), .Z(n3495) );
  MUX2_X1 U586 ( .A(n3798), .B(n530), .S(n560), .Z(n3494) );
  MUX2_X1 U587 ( .A(n3816), .B(n533), .S(n560), .Z(n3493) );
  MUX2_X1 U588 ( .A(n3834), .B(n536), .S(n560), .Z(n3492) );
  MUX2_X1 U589 ( .A(n3888), .B(n539), .S(n560), .Z(n3491) );
  MUX2_X1 U590 ( .A(n4086), .B(n542), .S(n560), .Z(n3490) );
  MUX2_X1 U591 ( .A(n4284), .B(n545), .S(n560), .Z(n3489) );
  OAI21_X1 U592 ( .B1(n872), .B2(n945), .A(n833), .ZN(n946) );
  MUX2_X1 U593 ( .A(n947), .B(n449), .S(n565), .Z(n3488) );
  MUX2_X1 U594 ( .A(n949), .B(n455), .S(n565), .Z(n3487) );
  MUX2_X1 U595 ( .A(n950), .B(n458), .S(n565), .Z(n3486) );
  MUX2_X1 U596 ( .A(n951), .B(n461), .S(n565), .Z(n3485) );
  MUX2_X1 U597 ( .A(n952), .B(n464), .S(n565), .Z(n3484) );
  MUX2_X1 U598 ( .A(n953), .B(n467), .S(n565), .Z(n3483) );
  MUX2_X1 U599 ( .A(n954), .B(n470), .S(n565), .Z(n3482) );
  MUX2_X1 U600 ( .A(n955), .B(n473), .S(n565), .Z(n3481) );
  MUX2_X1 U601 ( .A(n956), .B(n476), .S(n564), .Z(n3480) );
  MUX2_X1 U602 ( .A(n957), .B(n479), .S(n564), .Z(n3479) );
  MUX2_X1 U603 ( .A(n958), .B(n482), .S(n564), .Z(n3478) );
  MUX2_X1 U604 ( .A(n959), .B(n485), .S(n564), .Z(n3477) );
  MUX2_X1 U605 ( .A(n960), .B(n488), .S(n564), .Z(n3476) );
  MUX2_X1 U606 ( .A(n961), .B(n491), .S(n564), .Z(n3475) );
  MUX2_X1 U607 ( .A(n962), .B(n494), .S(n564), .Z(n3474) );
  MUX2_X1 U608 ( .A(n963), .B(n497), .S(n564), .Z(n3473) );
  MUX2_X1 U609 ( .A(n964), .B(n500), .S(n564), .Z(n3472) );
  MUX2_X1 U610 ( .A(n965), .B(n503), .S(n564), .Z(n3471) );
  MUX2_X1 U611 ( .A(n966), .B(n506), .S(n564), .Z(n3470) );
  MUX2_X1 U612 ( .A(n967), .B(n509), .S(n564), .Z(n3469) );
  MUX2_X1 U613 ( .A(n968), .B(n512), .S(n563), .Z(n3468) );
  MUX2_X1 U614 ( .A(n969), .B(n515), .S(n563), .Z(n3467) );
  MUX2_X1 U615 ( .A(n970), .B(n518), .S(n563), .Z(n3466) );
  MUX2_X1 U616 ( .A(n971), .B(n521), .S(n563), .Z(n3465) );
  MUX2_X1 U617 ( .A(n972), .B(n524), .S(n563), .Z(n3464) );
  MUX2_X1 U618 ( .A(n973), .B(n527), .S(n563), .Z(n3463) );
  MUX2_X1 U619 ( .A(n974), .B(n530), .S(n563), .Z(n3462) );
  MUX2_X1 U620 ( .A(n975), .B(n533), .S(n563), .Z(n3461) );
  MUX2_X1 U621 ( .A(n976), .B(n536), .S(n563), .Z(n3460) );
  MUX2_X1 U622 ( .A(n977), .B(n539), .S(n563), .Z(n3459) );
  MUX2_X1 U623 ( .A(n978), .B(n542), .S(n563), .Z(n3458) );
  MUX2_X1 U624 ( .A(n979), .B(n545), .S(n563), .Z(n3457) );
  OAI21_X1 U625 ( .B1(n906), .B2(n945), .A(n833), .ZN(n948) );
  MUX2_X1 U626 ( .A(n980), .B(n449), .S(n568), .Z(n3456) );
  MUX2_X1 U627 ( .A(n982), .B(n455), .S(n568), .Z(n3455) );
  MUX2_X1 U628 ( .A(n983), .B(n458), .S(n568), .Z(n3454) );
  MUX2_X1 U629 ( .A(n984), .B(n461), .S(n568), .Z(n3453) );
  MUX2_X1 U630 ( .A(n985), .B(n464), .S(n568), .Z(n3452) );
  MUX2_X1 U631 ( .A(n986), .B(n467), .S(n568), .Z(n3451) );
  MUX2_X1 U632 ( .A(n987), .B(n470), .S(n568), .Z(n3450) );
  MUX2_X1 U633 ( .A(n988), .B(n473), .S(n568), .Z(n3449) );
  MUX2_X1 U634 ( .A(n989), .B(n476), .S(n567), .Z(n3448) );
  MUX2_X1 U635 ( .A(n990), .B(n479), .S(n567), .Z(n3447) );
  MUX2_X1 U636 ( .A(n991), .B(n482), .S(n567), .Z(n3446) );
  MUX2_X1 U637 ( .A(n992), .B(n485), .S(n567), .Z(n3445) );
  MUX2_X1 U638 ( .A(n993), .B(n488), .S(n567), .Z(n3444) );
  MUX2_X1 U639 ( .A(n994), .B(n491), .S(n567), .Z(n3443) );
  MUX2_X1 U640 ( .A(n995), .B(n494), .S(n567), .Z(n3442) );
  MUX2_X1 U641 ( .A(n996), .B(n497), .S(n567), .Z(n3441) );
  MUX2_X1 U642 ( .A(n997), .B(n500), .S(n567), .Z(n3440) );
  MUX2_X1 U643 ( .A(n998), .B(n503), .S(n567), .Z(n3439) );
  MUX2_X1 U644 ( .A(n999), .B(n506), .S(n567), .Z(n3438) );
  MUX2_X1 U645 ( .A(n1000), .B(n509), .S(n567), .Z(n3437) );
  MUX2_X1 U646 ( .A(n1001), .B(n512), .S(n566), .Z(n3436) );
  MUX2_X1 U647 ( .A(n1002), .B(n515), .S(n566), .Z(n3435) );
  MUX2_X1 U648 ( .A(n1003), .B(n518), .S(n566), .Z(n3434) );
  MUX2_X1 U649 ( .A(n1004), .B(n521), .S(n566), .Z(n3433) );
  MUX2_X1 U650 ( .A(n1005), .B(n524), .S(n566), .Z(n3432) );
  MUX2_X1 U651 ( .A(n1006), .B(n527), .S(n566), .Z(n3431) );
  MUX2_X1 U652 ( .A(n1007), .B(n530), .S(n566), .Z(n3430) );
  MUX2_X1 U653 ( .A(n1008), .B(n533), .S(n566), .Z(n3429) );
  MUX2_X1 U654 ( .A(n1009), .B(n536), .S(n566), .Z(n3428) );
  MUX2_X1 U655 ( .A(n1010), .B(n539), .S(n566), .Z(n3427) );
  MUX2_X1 U656 ( .A(n1011), .B(n542), .S(n566), .Z(n3426) );
  MUX2_X1 U657 ( .A(n1012), .B(n545), .S(n566), .Z(n3425) );
  OAI21_X1 U658 ( .B1(n940), .B2(n945), .A(n833), .ZN(n981) );
  NAND3_X1 U659 ( .A1(n943), .A2(n942), .A3(ADD_WR[2]), .ZN(n945) );
  MUX2_X1 U660 ( .A(n3851), .B(n449), .S(n571), .Z(n3424) );
  MUX2_X1 U661 ( .A(n3869), .B(n455), .S(n571), .Z(n3423) );
  MUX2_X1 U662 ( .A(n3905), .B(n458), .S(n571), .Z(n3422) );
  MUX2_X1 U663 ( .A(n3923), .B(n461), .S(n571), .Z(n3421) );
  MUX2_X1 U664 ( .A(n3941), .B(n464), .S(n571), .Z(n3420) );
  MUX2_X1 U665 ( .A(n3959), .B(n467), .S(n571), .Z(n3419) );
  MUX2_X1 U666 ( .A(n3977), .B(n470), .S(n571), .Z(n3418) );
  MUX2_X1 U667 ( .A(n3995), .B(n473), .S(n571), .Z(n3417) );
  MUX2_X1 U668 ( .A(n4013), .B(n476), .S(n570), .Z(n3416) );
  MUX2_X1 U669 ( .A(n4031), .B(n479), .S(n570), .Z(n3415) );
  MUX2_X1 U670 ( .A(n4049), .B(n482), .S(n570), .Z(n3414) );
  MUX2_X1 U671 ( .A(n4067), .B(n485), .S(n570), .Z(n3413) );
  MUX2_X1 U672 ( .A(n4103), .B(n488), .S(n570), .Z(n3412) );
  MUX2_X1 U673 ( .A(n4121), .B(n491), .S(n570), .Z(n3411) );
  MUX2_X1 U674 ( .A(n4139), .B(n494), .S(n570), .Z(n3410) );
  MUX2_X1 U675 ( .A(n4157), .B(n497), .S(n570), .Z(n3409) );
  MUX2_X1 U676 ( .A(n4175), .B(n500), .S(n570), .Z(n3408) );
  MUX2_X1 U677 ( .A(n4193), .B(n503), .S(n570), .Z(n3407) );
  MUX2_X1 U678 ( .A(n4211), .B(n506), .S(n570), .Z(n3406) );
  MUX2_X1 U679 ( .A(n4229), .B(n509), .S(n570), .Z(n3405) );
  MUX2_X1 U680 ( .A(n4247), .B(n512), .S(n569), .Z(n3404) );
  MUX2_X1 U681 ( .A(n4265), .B(n515), .S(n569), .Z(n3403) );
  MUX2_X1 U682 ( .A(n3725), .B(n518), .S(n569), .Z(n3402) );
  MUX2_X1 U683 ( .A(n3743), .B(n521), .S(n569), .Z(n3401) );
  MUX2_X1 U684 ( .A(n3761), .B(n524), .S(n569), .Z(n3400) );
  MUX2_X1 U685 ( .A(n3779), .B(n527), .S(n569), .Z(n3399) );
  MUX2_X1 U686 ( .A(n3797), .B(n530), .S(n569), .Z(n3398) );
  MUX2_X1 U687 ( .A(n3815), .B(n533), .S(n569), .Z(n3397) );
  MUX2_X1 U688 ( .A(n3833), .B(n536), .S(n569), .Z(n3396) );
  MUX2_X1 U689 ( .A(n3887), .B(n539), .S(n569), .Z(n3395) );
  MUX2_X1 U690 ( .A(n4085), .B(n542), .S(n569), .Z(n3394) );
  MUX2_X1 U691 ( .A(n4283), .B(n545), .S(n569), .Z(n3393) );
  OAI21_X1 U692 ( .B1(n870), .B2(n1014), .A(n833), .ZN(n1013) );
  MUX2_X1 U693 ( .A(n3850), .B(n449), .S(n574), .Z(n3392) );
  MUX2_X1 U694 ( .A(n3868), .B(n455), .S(n574), .Z(n3391) );
  MUX2_X1 U695 ( .A(n3904), .B(n458), .S(n574), .Z(n3390) );
  MUX2_X1 U696 ( .A(n3922), .B(n461), .S(n574), .Z(n3389) );
  MUX2_X1 U697 ( .A(n3940), .B(n464), .S(n574), .Z(n3388) );
  MUX2_X1 U698 ( .A(n3958), .B(n467), .S(n574), .Z(n3387) );
  MUX2_X1 U699 ( .A(n3976), .B(n470), .S(n574), .Z(n3386) );
  MUX2_X1 U700 ( .A(n3994), .B(n473), .S(n574), .Z(n3385) );
  MUX2_X1 U701 ( .A(n4012), .B(n476), .S(n573), .Z(n3384) );
  MUX2_X1 U702 ( .A(n4030), .B(n479), .S(n573), .Z(n3383) );
  MUX2_X1 U703 ( .A(n4048), .B(n482), .S(n573), .Z(n3382) );
  MUX2_X1 U704 ( .A(n4066), .B(n485), .S(n573), .Z(n3381) );
  MUX2_X1 U705 ( .A(n4102), .B(n488), .S(n573), .Z(n3380) );
  MUX2_X1 U706 ( .A(n4120), .B(n491), .S(n573), .Z(n3379) );
  MUX2_X1 U707 ( .A(n4138), .B(n494), .S(n573), .Z(n3378) );
  MUX2_X1 U708 ( .A(n4156), .B(n497), .S(n573), .Z(n3377) );
  MUX2_X1 U709 ( .A(n4174), .B(n500), .S(n573), .Z(n3376) );
  MUX2_X1 U710 ( .A(n4192), .B(n503), .S(n573), .Z(n3375) );
  MUX2_X1 U711 ( .A(n4210), .B(n506), .S(n573), .Z(n3374) );
  MUX2_X1 U712 ( .A(n4228), .B(n509), .S(n573), .Z(n3373) );
  MUX2_X1 U713 ( .A(n4246), .B(n512), .S(n572), .Z(n3372) );
  MUX2_X1 U714 ( .A(n4264), .B(n515), .S(n572), .Z(n3371) );
  MUX2_X1 U715 ( .A(n3724), .B(n518), .S(n572), .Z(n3370) );
  MUX2_X1 U716 ( .A(n3742), .B(n521), .S(n572), .Z(n3369) );
  MUX2_X1 U717 ( .A(n3760), .B(n524), .S(n572), .Z(n3368) );
  MUX2_X1 U718 ( .A(n3778), .B(n527), .S(n572), .Z(n3367) );
  MUX2_X1 U719 ( .A(n3796), .B(n530), .S(n572), .Z(n3366) );
  MUX2_X1 U720 ( .A(n3814), .B(n533), .S(n572), .Z(n3365) );
  MUX2_X1 U721 ( .A(n3832), .B(n536), .S(n572), .Z(n3364) );
  MUX2_X1 U722 ( .A(n3886), .B(n539), .S(n572), .Z(n3363) );
  MUX2_X1 U723 ( .A(n4084), .B(n542), .S(n572), .Z(n3362) );
  MUX2_X1 U724 ( .A(n4282), .B(n545), .S(n572), .Z(n3361) );
  OAI21_X1 U725 ( .B1(n872), .B2(n1014), .A(n833), .ZN(n1015) );
  MUX2_X1 U726 ( .A(n1016), .B(n449), .S(n577), .Z(n3360) );
  MUX2_X1 U727 ( .A(n1018), .B(n455), .S(n577), .Z(n3359) );
  MUX2_X1 U728 ( .A(n1019), .B(n458), .S(n577), .Z(n3358) );
  MUX2_X1 U729 ( .A(n1020), .B(n461), .S(n577), .Z(n3357) );
  MUX2_X1 U730 ( .A(n1021), .B(n464), .S(n577), .Z(n3356) );
  MUX2_X1 U731 ( .A(n1022), .B(n467), .S(n577), .Z(n3355) );
  MUX2_X1 U732 ( .A(n1023), .B(n470), .S(n577), .Z(n3354) );
  MUX2_X1 U733 ( .A(n1024), .B(n473), .S(n577), .Z(n3353) );
  MUX2_X1 U734 ( .A(n1025), .B(n476), .S(n576), .Z(n3352) );
  MUX2_X1 U735 ( .A(n1026), .B(n479), .S(n576), .Z(n3351) );
  MUX2_X1 U736 ( .A(n1027), .B(n482), .S(n576), .Z(n3350) );
  MUX2_X1 U737 ( .A(n1028), .B(n485), .S(n576), .Z(n3349) );
  MUX2_X1 U738 ( .A(n1029), .B(n488), .S(n576), .Z(n3348) );
  MUX2_X1 U739 ( .A(n1030), .B(n491), .S(n576), .Z(n3347) );
  MUX2_X1 U740 ( .A(n1031), .B(n494), .S(n576), .Z(n3346) );
  MUX2_X1 U741 ( .A(n1032), .B(n497), .S(n576), .Z(n3345) );
  MUX2_X1 U742 ( .A(n1033), .B(n500), .S(n576), .Z(n3344) );
  MUX2_X1 U743 ( .A(n1034), .B(n503), .S(n576), .Z(n3343) );
  MUX2_X1 U744 ( .A(n1035), .B(n506), .S(n576), .Z(n3342) );
  MUX2_X1 U745 ( .A(n1036), .B(n509), .S(n576), .Z(n3341) );
  MUX2_X1 U746 ( .A(n1037), .B(n512), .S(n575), .Z(n3340) );
  MUX2_X1 U747 ( .A(n1038), .B(n515), .S(n575), .Z(n3339) );
  MUX2_X1 U748 ( .A(n1039), .B(n518), .S(n575), .Z(n3338) );
  MUX2_X1 U749 ( .A(n1040), .B(n521), .S(n575), .Z(n3337) );
  MUX2_X1 U750 ( .A(n1041), .B(n524), .S(n575), .Z(n3336) );
  MUX2_X1 U751 ( .A(n1042), .B(n527), .S(n575), .Z(n3335) );
  MUX2_X1 U752 ( .A(n1043), .B(n530), .S(n575), .Z(n3334) );
  MUX2_X1 U753 ( .A(n1044), .B(n533), .S(n575), .Z(n3333) );
  MUX2_X1 U754 ( .A(n1045), .B(n536), .S(n575), .Z(n3332) );
  MUX2_X1 U755 ( .A(n1046), .B(n539), .S(n575), .Z(n3331) );
  MUX2_X1 U756 ( .A(n1047), .B(n542), .S(n575), .Z(n3330) );
  MUX2_X1 U757 ( .A(n1048), .B(n545), .S(n575), .Z(n3329) );
  OAI21_X1 U758 ( .B1(n906), .B2(n1014), .A(n833), .ZN(n1017) );
  MUX2_X1 U759 ( .A(n1049), .B(n450), .S(n580), .Z(n3328) );
  MUX2_X1 U760 ( .A(n1051), .B(n456), .S(n580), .Z(n3327) );
  MUX2_X1 U761 ( .A(n1052), .B(n459), .S(n580), .Z(n3326) );
  MUX2_X1 U762 ( .A(n1053), .B(n462), .S(n580), .Z(n3325) );
  MUX2_X1 U763 ( .A(n1054), .B(n465), .S(n580), .Z(n3324) );
  MUX2_X1 U764 ( .A(n1055), .B(n468), .S(n580), .Z(n3323) );
  MUX2_X1 U765 ( .A(n1056), .B(n471), .S(n580), .Z(n3322) );
  MUX2_X1 U766 ( .A(n1057), .B(n474), .S(n580), .Z(n3321) );
  MUX2_X1 U767 ( .A(n1058), .B(n477), .S(n579), .Z(n3320) );
  MUX2_X1 U768 ( .A(n1059), .B(n480), .S(n579), .Z(n3319) );
  MUX2_X1 U769 ( .A(n1060), .B(n483), .S(n579), .Z(n3318) );
  MUX2_X1 U770 ( .A(n1061), .B(n486), .S(n579), .Z(n3317) );
  MUX2_X1 U771 ( .A(n1062), .B(n489), .S(n579), .Z(n3316) );
  MUX2_X1 U772 ( .A(n1063), .B(n492), .S(n579), .Z(n3315) );
  MUX2_X1 U773 ( .A(n1064), .B(n495), .S(n579), .Z(n3314) );
  MUX2_X1 U774 ( .A(n1065), .B(n498), .S(n579), .Z(n3313) );
  MUX2_X1 U775 ( .A(n1066), .B(n501), .S(n579), .Z(n3312) );
  MUX2_X1 U776 ( .A(n1067), .B(n504), .S(n579), .Z(n3311) );
  MUX2_X1 U777 ( .A(n1068), .B(n507), .S(n579), .Z(n3310) );
  MUX2_X1 U778 ( .A(n1069), .B(n510), .S(n579), .Z(n3309) );
  MUX2_X1 U779 ( .A(n1070), .B(n513), .S(n578), .Z(n3308) );
  MUX2_X1 U780 ( .A(n1071), .B(n516), .S(n578), .Z(n3307) );
  MUX2_X1 U781 ( .A(n1072), .B(n519), .S(n578), .Z(n3306) );
  MUX2_X1 U782 ( .A(n1073), .B(n522), .S(n578), .Z(n3305) );
  MUX2_X1 U783 ( .A(n1074), .B(n525), .S(n578), .Z(n3304) );
  MUX2_X1 U784 ( .A(n1075), .B(n528), .S(n578), .Z(n3303) );
  MUX2_X1 U785 ( .A(n1076), .B(n531), .S(n578), .Z(n3302) );
  MUX2_X1 U786 ( .A(n1077), .B(n534), .S(n578), .Z(n3301) );
  MUX2_X1 U787 ( .A(n1078), .B(n537), .S(n578), .Z(n3300) );
  MUX2_X1 U788 ( .A(n1079), .B(n540), .S(n578), .Z(n3299) );
  MUX2_X1 U789 ( .A(n1080), .B(n543), .S(n578), .Z(n3298) );
  MUX2_X1 U790 ( .A(n1081), .B(n546), .S(n578), .Z(n3297) );
  OAI21_X1 U791 ( .B1(n940), .B2(n1014), .A(n833), .ZN(n1050) );
  NAND3_X1 U792 ( .A1(n943), .A2(n941), .A3(ADD_WR[3]), .ZN(n1014) );
  MUX2_X1 U793 ( .A(n3849), .B(n450), .S(n583), .Z(n3296) );
  MUX2_X1 U794 ( .A(n3867), .B(n456), .S(n583), .Z(n3295) );
  MUX2_X1 U795 ( .A(n3903), .B(n459), .S(n583), .Z(n3294) );
  MUX2_X1 U796 ( .A(n3921), .B(n462), .S(n583), .Z(n3293) );
  MUX2_X1 U797 ( .A(n3939), .B(n465), .S(n583), .Z(n3292) );
  MUX2_X1 U798 ( .A(n3957), .B(n468), .S(n583), .Z(n3291) );
  MUX2_X1 U799 ( .A(n3975), .B(n471), .S(n583), .Z(n3290) );
  MUX2_X1 U800 ( .A(n3993), .B(n474), .S(n583), .Z(n3289) );
  MUX2_X1 U801 ( .A(n4011), .B(n477), .S(n582), .Z(n3288) );
  MUX2_X1 U802 ( .A(n4029), .B(n480), .S(n582), .Z(n3287) );
  MUX2_X1 U803 ( .A(n4047), .B(n483), .S(n582), .Z(n3286) );
  MUX2_X1 U804 ( .A(n4065), .B(n486), .S(n582), .Z(n3285) );
  MUX2_X1 U805 ( .A(n4101), .B(n489), .S(n582), .Z(n3284) );
  MUX2_X1 U806 ( .A(n4119), .B(n492), .S(n582), .Z(n3283) );
  MUX2_X1 U807 ( .A(n4137), .B(n495), .S(n582), .Z(n3282) );
  MUX2_X1 U808 ( .A(n4155), .B(n498), .S(n582), .Z(n3281) );
  MUX2_X1 U809 ( .A(n4173), .B(n501), .S(n582), .Z(n3280) );
  MUX2_X1 U810 ( .A(n4191), .B(n504), .S(n582), .Z(n3279) );
  MUX2_X1 U811 ( .A(n4209), .B(n507), .S(n582), .Z(n3278) );
  MUX2_X1 U812 ( .A(n4227), .B(n510), .S(n582), .Z(n3277) );
  MUX2_X1 U813 ( .A(n4245), .B(n513), .S(n581), .Z(n3276) );
  MUX2_X1 U814 ( .A(n4263), .B(n516), .S(n581), .Z(n3275) );
  MUX2_X1 U815 ( .A(n3723), .B(n519), .S(n581), .Z(n3274) );
  MUX2_X1 U816 ( .A(n3741), .B(n522), .S(n581), .Z(n3273) );
  MUX2_X1 U817 ( .A(n3759), .B(n525), .S(n581), .Z(n3272) );
  MUX2_X1 U818 ( .A(n3777), .B(n528), .S(n581), .Z(n3271) );
  MUX2_X1 U819 ( .A(n3795), .B(n531), .S(n581), .Z(n3270) );
  MUX2_X1 U820 ( .A(n3813), .B(n534), .S(n581), .Z(n3269) );
  MUX2_X1 U821 ( .A(n3831), .B(n537), .S(n581), .Z(n3268) );
  MUX2_X1 U822 ( .A(n3885), .B(n540), .S(n581), .Z(n3267) );
  MUX2_X1 U823 ( .A(n4083), .B(n543), .S(n581), .Z(n3266) );
  MUX2_X1 U824 ( .A(n4281), .B(n546), .S(n581), .Z(n3265) );
  OAI21_X1 U825 ( .B1(n870), .B2(n1083), .A(n833), .ZN(n1082) );
  MUX2_X1 U826 ( .A(n3848), .B(n450), .S(n586), .Z(n3264) );
  MUX2_X1 U827 ( .A(n3866), .B(n456), .S(n586), .Z(n3263) );
  MUX2_X1 U828 ( .A(n3902), .B(n459), .S(n586), .Z(n3262) );
  MUX2_X1 U829 ( .A(n3920), .B(n462), .S(n586), .Z(n3261) );
  MUX2_X1 U830 ( .A(n3938), .B(n465), .S(n586), .Z(n3260) );
  MUX2_X1 U831 ( .A(n3956), .B(n468), .S(n586), .Z(n3259) );
  MUX2_X1 U832 ( .A(n3974), .B(n471), .S(n586), .Z(n3258) );
  MUX2_X1 U833 ( .A(n3992), .B(n474), .S(n586), .Z(n3257) );
  MUX2_X1 U834 ( .A(n4010), .B(n477), .S(n585), .Z(n3256) );
  MUX2_X1 U835 ( .A(n4028), .B(n480), .S(n585), .Z(n3255) );
  MUX2_X1 U836 ( .A(n4046), .B(n483), .S(n585), .Z(n3254) );
  MUX2_X1 U837 ( .A(n4064), .B(n486), .S(n585), .Z(n3253) );
  MUX2_X1 U838 ( .A(n4100), .B(n489), .S(n585), .Z(n3252) );
  MUX2_X1 U839 ( .A(n4118), .B(n492), .S(n585), .Z(n3251) );
  MUX2_X1 U840 ( .A(n4136), .B(n495), .S(n585), .Z(n3250) );
  MUX2_X1 U841 ( .A(n4154), .B(n498), .S(n585), .Z(n3249) );
  MUX2_X1 U842 ( .A(n4172), .B(n501), .S(n585), .Z(n3248) );
  MUX2_X1 U843 ( .A(n4190), .B(n504), .S(n585), .Z(n3247) );
  MUX2_X1 U844 ( .A(n4208), .B(n507), .S(n585), .Z(n3246) );
  MUX2_X1 U845 ( .A(n4226), .B(n510), .S(n585), .Z(n3245) );
  MUX2_X1 U846 ( .A(n4244), .B(n513), .S(n584), .Z(n3244) );
  MUX2_X1 U847 ( .A(n4262), .B(n516), .S(n584), .Z(n3243) );
  MUX2_X1 U848 ( .A(n3722), .B(n519), .S(n584), .Z(n3242) );
  MUX2_X1 U849 ( .A(n3740), .B(n522), .S(n584), .Z(n3241) );
  MUX2_X1 U850 ( .A(n3758), .B(n525), .S(n584), .Z(n3240) );
  MUX2_X1 U851 ( .A(n3776), .B(n528), .S(n584), .Z(n3239) );
  MUX2_X1 U852 ( .A(n3794), .B(n531), .S(n584), .Z(n3238) );
  MUX2_X1 U853 ( .A(n3812), .B(n534), .S(n584), .Z(n3237) );
  MUX2_X1 U854 ( .A(n3830), .B(n537), .S(n584), .Z(n3236) );
  MUX2_X1 U855 ( .A(n3884), .B(n540), .S(n584), .Z(n3235) );
  MUX2_X1 U856 ( .A(n4082), .B(n543), .S(n584), .Z(n3234) );
  MUX2_X1 U857 ( .A(n4280), .B(n546), .S(n584), .Z(n3233) );
  OAI21_X1 U858 ( .B1(n872), .B2(n1083), .A(RESET), .ZN(n1084) );
  MUX2_X1 U859 ( .A(n1085), .B(n450), .S(n589), .Z(n3232) );
  MUX2_X1 U860 ( .A(n1087), .B(n456), .S(n589), .Z(n3231) );
  MUX2_X1 U861 ( .A(n1088), .B(n459), .S(n589), .Z(n3230) );
  MUX2_X1 U862 ( .A(n1089), .B(n462), .S(n589), .Z(n3229) );
  MUX2_X1 U863 ( .A(n1090), .B(n465), .S(n589), .Z(n3228) );
  MUX2_X1 U864 ( .A(n1091), .B(n468), .S(n589), .Z(n3227) );
  MUX2_X1 U865 ( .A(n1092), .B(n471), .S(n589), .Z(n3226) );
  MUX2_X1 U866 ( .A(n1093), .B(n474), .S(n589), .Z(n3225) );
  MUX2_X1 U867 ( .A(n1094), .B(n477), .S(n588), .Z(n3224) );
  MUX2_X1 U868 ( .A(n1095), .B(n480), .S(n588), .Z(n3223) );
  MUX2_X1 U869 ( .A(n1096), .B(n483), .S(n588), .Z(n3222) );
  MUX2_X1 U870 ( .A(n1097), .B(n486), .S(n588), .Z(n3221) );
  MUX2_X1 U871 ( .A(n1098), .B(n489), .S(n588), .Z(n3220) );
  MUX2_X1 U872 ( .A(n1099), .B(n492), .S(n588), .Z(n3219) );
  MUX2_X1 U873 ( .A(n1100), .B(n495), .S(n588), .Z(n3218) );
  MUX2_X1 U874 ( .A(n1101), .B(n498), .S(n588), .Z(n3217) );
  MUX2_X1 U875 ( .A(n1102), .B(n501), .S(n588), .Z(n3216) );
  MUX2_X1 U876 ( .A(n1103), .B(n504), .S(n588), .Z(n3215) );
  MUX2_X1 U877 ( .A(n1104), .B(n507), .S(n588), .Z(n3214) );
  MUX2_X1 U878 ( .A(n1105), .B(n510), .S(n588), .Z(n3213) );
  MUX2_X1 U879 ( .A(n1106), .B(n513), .S(n587), .Z(n3212) );
  MUX2_X1 U880 ( .A(n1107), .B(n516), .S(n587), .Z(n3211) );
  MUX2_X1 U881 ( .A(n1108), .B(n519), .S(n587), .Z(n3210) );
  MUX2_X1 U882 ( .A(n1109), .B(n522), .S(n587), .Z(n3209) );
  MUX2_X1 U883 ( .A(n1110), .B(n525), .S(n587), .Z(n3208) );
  MUX2_X1 U884 ( .A(n1111), .B(n528), .S(n587), .Z(n3207) );
  MUX2_X1 U885 ( .A(n1112), .B(n531), .S(n587), .Z(n3206) );
  MUX2_X1 U886 ( .A(n1113), .B(n534), .S(n587), .Z(n3205) );
  MUX2_X1 U887 ( .A(n1114), .B(n537), .S(n587), .Z(n3204) );
  MUX2_X1 U888 ( .A(n1115), .B(n540), .S(n587), .Z(n3203) );
  MUX2_X1 U889 ( .A(n1116), .B(n543), .S(n587), .Z(n3202) );
  MUX2_X1 U890 ( .A(n1117), .B(n546), .S(n587), .Z(n3201) );
  OAI21_X1 U891 ( .B1(n906), .B2(n1083), .A(RESET), .ZN(n1086) );
  MUX2_X1 U892 ( .A(n1118), .B(n450), .S(n592), .Z(n3200) );
  MUX2_X1 U893 ( .A(n1120), .B(n456), .S(n592), .Z(n3199) );
  MUX2_X1 U894 ( .A(n1121), .B(n459), .S(n592), .Z(n3198) );
  MUX2_X1 U895 ( .A(n1122), .B(n462), .S(n592), .Z(n3197) );
  MUX2_X1 U896 ( .A(n1123), .B(n465), .S(n592), .Z(n3196) );
  MUX2_X1 U897 ( .A(n1124), .B(n468), .S(n592), .Z(n3195) );
  MUX2_X1 U898 ( .A(n1125), .B(n471), .S(n592), .Z(n3194) );
  MUX2_X1 U899 ( .A(n1126), .B(n474), .S(n592), .Z(n3193) );
  MUX2_X1 U900 ( .A(n1127), .B(n477), .S(n591), .Z(n3192) );
  MUX2_X1 U901 ( .A(n1128), .B(n480), .S(n591), .Z(n3191) );
  MUX2_X1 U902 ( .A(n1129), .B(n483), .S(n591), .Z(n3190) );
  MUX2_X1 U903 ( .A(n1130), .B(n486), .S(n591), .Z(n3189) );
  MUX2_X1 U904 ( .A(n1131), .B(n489), .S(n591), .Z(n3188) );
  MUX2_X1 U905 ( .A(n1132), .B(n492), .S(n591), .Z(n3187) );
  MUX2_X1 U906 ( .A(n1133), .B(n495), .S(n591), .Z(n3186) );
  MUX2_X1 U907 ( .A(n1134), .B(n498), .S(n591), .Z(n3185) );
  MUX2_X1 U908 ( .A(n1135), .B(n501), .S(n591), .Z(n3184) );
  MUX2_X1 U909 ( .A(n1136), .B(n504), .S(n591), .Z(n3183) );
  MUX2_X1 U910 ( .A(n1137), .B(n507), .S(n591), .Z(n3182) );
  MUX2_X1 U911 ( .A(n1138), .B(n510), .S(n591), .Z(n3181) );
  MUX2_X1 U912 ( .A(n1139), .B(n513), .S(n590), .Z(n3180) );
  MUX2_X1 U913 ( .A(n1140), .B(n516), .S(n590), .Z(n3179) );
  MUX2_X1 U914 ( .A(n1141), .B(n519), .S(n590), .Z(n3178) );
  MUX2_X1 U915 ( .A(n1142), .B(n522), .S(n590), .Z(n3177) );
  MUX2_X1 U916 ( .A(n1143), .B(n525), .S(n590), .Z(n3176) );
  MUX2_X1 U917 ( .A(n1144), .B(n528), .S(n590), .Z(n3175) );
  MUX2_X1 U918 ( .A(n1145), .B(n531), .S(n590), .Z(n3174) );
  MUX2_X1 U919 ( .A(n1146), .B(n534), .S(n590), .Z(n3173) );
  MUX2_X1 U920 ( .A(n1147), .B(n537), .S(n590), .Z(n3172) );
  MUX2_X1 U921 ( .A(n1148), .B(n540), .S(n590), .Z(n3171) );
  MUX2_X1 U922 ( .A(n1149), .B(n543), .S(n590), .Z(n3170) );
  MUX2_X1 U923 ( .A(n1150), .B(n546), .S(n590), .Z(n3169) );
  OAI21_X1 U924 ( .B1(n940), .B2(n1083), .A(RESET), .ZN(n1119) );
  NAND3_X1 U925 ( .A1(ADD_WR[2]), .A2(n943), .A3(ADD_WR[3]), .ZN(n1083) );
  NOR2_X1 U926 ( .A1(n1151), .A2(ADD_WR[4]), .ZN(n943) );
  MUX2_X1 U927 ( .A(n3858), .B(n450), .S(n595), .Z(n3168) );
  MUX2_X1 U928 ( .A(n3876), .B(n456), .S(n595), .Z(n3167) );
  MUX2_X1 U929 ( .A(n3912), .B(n459), .S(n595), .Z(n3166) );
  MUX2_X1 U930 ( .A(n3930), .B(n462), .S(n595), .Z(n3165) );
  MUX2_X1 U931 ( .A(n3948), .B(n465), .S(n595), .Z(n3164) );
  MUX2_X1 U932 ( .A(n3966), .B(n468), .S(n595), .Z(n3163) );
  MUX2_X1 U933 ( .A(n3984), .B(n471), .S(n595), .Z(n3162) );
  MUX2_X1 U934 ( .A(n4002), .B(n474), .S(n595), .Z(n3161) );
  MUX2_X1 U935 ( .A(n4020), .B(n477), .S(n594), .Z(n3160) );
  MUX2_X1 U936 ( .A(n4038), .B(n480), .S(n594), .Z(n3159) );
  MUX2_X1 U937 ( .A(n4056), .B(n483), .S(n594), .Z(n3158) );
  MUX2_X1 U938 ( .A(n4074), .B(n486), .S(n594), .Z(n3157) );
  MUX2_X1 U939 ( .A(n4110), .B(n489), .S(n594), .Z(n3156) );
  MUX2_X1 U940 ( .A(n4128), .B(n492), .S(n594), .Z(n3155) );
  MUX2_X1 U941 ( .A(n4146), .B(n495), .S(n594), .Z(n3154) );
  MUX2_X1 U942 ( .A(n4164), .B(n498), .S(n594), .Z(n3153) );
  MUX2_X1 U943 ( .A(n4182), .B(n501), .S(n594), .Z(n3152) );
  MUX2_X1 U944 ( .A(n4200), .B(n504), .S(n594), .Z(n3151) );
  MUX2_X1 U945 ( .A(n4218), .B(n507), .S(n594), .Z(n3150) );
  MUX2_X1 U946 ( .A(n4236), .B(n510), .S(n594), .Z(n3149) );
  MUX2_X1 U947 ( .A(n4254), .B(n513), .S(n593), .Z(n3148) );
  MUX2_X1 U948 ( .A(n4272), .B(n516), .S(n593), .Z(n3147) );
  MUX2_X1 U949 ( .A(n3732), .B(n519), .S(n593), .Z(n3146) );
  MUX2_X1 U950 ( .A(n3750), .B(n522), .S(n593), .Z(n3145) );
  MUX2_X1 U951 ( .A(n3768), .B(n525), .S(n593), .Z(n3144) );
  MUX2_X1 U952 ( .A(n3786), .B(n528), .S(n593), .Z(n3143) );
  MUX2_X1 U953 ( .A(n3804), .B(n531), .S(n593), .Z(n3142) );
  MUX2_X1 U954 ( .A(n3822), .B(n534), .S(n593), .Z(n3141) );
  MUX2_X1 U955 ( .A(n3840), .B(n537), .S(n593), .Z(n3140) );
  MUX2_X1 U956 ( .A(n3894), .B(n540), .S(n593), .Z(n3139) );
  MUX2_X1 U957 ( .A(n4092), .B(n543), .S(n593), .Z(n3138) );
  MUX2_X1 U958 ( .A(n4290), .B(n546), .S(n593), .Z(n3137) );
  OAI21_X1 U959 ( .B1(n870), .B2(n1153), .A(n833), .ZN(n1152) );
  MUX2_X1 U960 ( .A(n3859), .B(n450), .S(n598), .Z(n3136) );
  MUX2_X1 U961 ( .A(n3877), .B(n456), .S(n598), .Z(n3135) );
  MUX2_X1 U962 ( .A(n3913), .B(n459), .S(n598), .Z(n3134) );
  MUX2_X1 U963 ( .A(n3931), .B(n462), .S(n598), .Z(n3133) );
  MUX2_X1 U964 ( .A(n3949), .B(n465), .S(n598), .Z(n3132) );
  MUX2_X1 U965 ( .A(n3967), .B(n468), .S(n598), .Z(n3131) );
  MUX2_X1 U966 ( .A(n3985), .B(n471), .S(n598), .Z(n3130) );
  MUX2_X1 U967 ( .A(n4003), .B(n474), .S(n598), .Z(n3129) );
  MUX2_X1 U968 ( .A(n4021), .B(n477), .S(n597), .Z(n3128) );
  MUX2_X1 U969 ( .A(n4039), .B(n480), .S(n597), .Z(n3127) );
  MUX2_X1 U970 ( .A(n4057), .B(n483), .S(n597), .Z(n3126) );
  MUX2_X1 U971 ( .A(n4075), .B(n486), .S(n597), .Z(n3125) );
  MUX2_X1 U972 ( .A(n4111), .B(n489), .S(n597), .Z(n3124) );
  MUX2_X1 U973 ( .A(n4129), .B(n492), .S(n597), .Z(n3123) );
  MUX2_X1 U974 ( .A(n4147), .B(n495), .S(n597), .Z(n3122) );
  MUX2_X1 U975 ( .A(n4165), .B(n498), .S(n597), .Z(n3121) );
  MUX2_X1 U976 ( .A(n4183), .B(n501), .S(n597), .Z(n3120) );
  MUX2_X1 U977 ( .A(n4201), .B(n504), .S(n597), .Z(n3119) );
  MUX2_X1 U978 ( .A(n4219), .B(n507), .S(n597), .Z(n3118) );
  MUX2_X1 U979 ( .A(n4237), .B(n510), .S(n597), .Z(n3117) );
  MUX2_X1 U980 ( .A(n4255), .B(n513), .S(n596), .Z(n3116) );
  MUX2_X1 U981 ( .A(n4273), .B(n516), .S(n596), .Z(n3115) );
  MUX2_X1 U982 ( .A(n3733), .B(n519), .S(n596), .Z(n3114) );
  MUX2_X1 U983 ( .A(n3751), .B(n522), .S(n596), .Z(n3113) );
  MUX2_X1 U984 ( .A(n3769), .B(n525), .S(n596), .Z(n3112) );
  MUX2_X1 U985 ( .A(n3787), .B(n528), .S(n596), .Z(n3111) );
  MUX2_X1 U986 ( .A(n3805), .B(n531), .S(n596), .Z(n3110) );
  MUX2_X1 U987 ( .A(n3823), .B(n534), .S(n596), .Z(n3109) );
  MUX2_X1 U988 ( .A(n3841), .B(n537), .S(n596), .Z(n3108) );
  MUX2_X1 U989 ( .A(n3895), .B(n540), .S(n596), .Z(n3107) );
  MUX2_X1 U990 ( .A(n4093), .B(n543), .S(n596), .Z(n3106) );
  MUX2_X1 U991 ( .A(n4291), .B(n546), .S(n596), .Z(n3105) );
  OAI21_X1 U992 ( .B1(n872), .B2(n1153), .A(RESET), .ZN(n1154) );
  MUX2_X1 U993 ( .A(n1155), .B(n450), .S(n601), .Z(n3104) );
  MUX2_X1 U994 ( .A(n1157), .B(n456), .S(n601), .Z(n3103) );
  MUX2_X1 U995 ( .A(n1158), .B(n459), .S(n601), .Z(n3102) );
  MUX2_X1 U996 ( .A(n1159), .B(n462), .S(n601), .Z(n3101) );
  MUX2_X1 U997 ( .A(n1160), .B(n465), .S(n601), .Z(n3100) );
  MUX2_X1 U998 ( .A(n1161), .B(n468), .S(n601), .Z(n3099) );
  MUX2_X1 U999 ( .A(n1162), .B(n471), .S(n601), .Z(n3098) );
  MUX2_X1 U1000 ( .A(n1163), .B(n474), .S(n601), .Z(n3097) );
  MUX2_X1 U1001 ( .A(n1164), .B(n477), .S(n600), .Z(n3096) );
  MUX2_X1 U1002 ( .A(n1165), .B(n480), .S(n600), .Z(n3095) );
  MUX2_X1 U1003 ( .A(n1166), .B(n483), .S(n600), .Z(n3094) );
  MUX2_X1 U1004 ( .A(n1167), .B(n486), .S(n600), .Z(n3093) );
  MUX2_X1 U1005 ( .A(n1168), .B(n489), .S(n600), .Z(n3092) );
  MUX2_X1 U1006 ( .A(n1169), .B(n492), .S(n600), .Z(n3091) );
  MUX2_X1 U1007 ( .A(n1170), .B(n495), .S(n600), .Z(n3090) );
  MUX2_X1 U1008 ( .A(n1171), .B(n498), .S(n600), .Z(n3089) );
  MUX2_X1 U1009 ( .A(n1172), .B(n501), .S(n600), .Z(n3088) );
  MUX2_X1 U1010 ( .A(n1173), .B(n504), .S(n600), .Z(n3087) );
  MUX2_X1 U1011 ( .A(n1174), .B(n507), .S(n600), .Z(n3086) );
  MUX2_X1 U1012 ( .A(n1175), .B(n510), .S(n600), .Z(n3085) );
  MUX2_X1 U1013 ( .A(n1176), .B(n513), .S(n599), .Z(n3084) );
  MUX2_X1 U1014 ( .A(n1177), .B(n516), .S(n599), .Z(n3083) );
  MUX2_X1 U1015 ( .A(n1178), .B(n519), .S(n599), .Z(n3082) );
  MUX2_X1 U1016 ( .A(n1179), .B(n522), .S(n599), .Z(n3081) );
  MUX2_X1 U1017 ( .A(n1180), .B(n525), .S(n599), .Z(n3080) );
  MUX2_X1 U1018 ( .A(n1181), .B(n528), .S(n599), .Z(n3079) );
  MUX2_X1 U1019 ( .A(n1182), .B(n531), .S(n599), .Z(n3078) );
  MUX2_X1 U1020 ( .A(n1183), .B(n534), .S(n599), .Z(n3077) );
  MUX2_X1 U1021 ( .A(n1184), .B(n537), .S(n599), .Z(n3076) );
  MUX2_X1 U1022 ( .A(n1185), .B(n540), .S(n599), .Z(n3075) );
  MUX2_X1 U1023 ( .A(n1186), .B(n543), .S(n599), .Z(n3074) );
  MUX2_X1 U1024 ( .A(n1187), .B(n546), .S(n599), .Z(n3073) );
  OAI21_X1 U1025 ( .B1(n906), .B2(n1153), .A(RESET), .ZN(n1156) );
  MUX2_X1 U1026 ( .A(n1188), .B(n450), .S(n604), .Z(n3072) );
  MUX2_X1 U1027 ( .A(n1190), .B(n456), .S(n604), .Z(n3071) );
  MUX2_X1 U1028 ( .A(n1191), .B(n459), .S(n604), .Z(n3070) );
  MUX2_X1 U1029 ( .A(n1192), .B(n462), .S(n604), .Z(n3069) );
  MUX2_X1 U1030 ( .A(n1193), .B(n465), .S(n604), .Z(n3068) );
  MUX2_X1 U1031 ( .A(n1194), .B(n468), .S(n604), .Z(n3067) );
  MUX2_X1 U1032 ( .A(n1195), .B(n471), .S(n604), .Z(n3066) );
  MUX2_X1 U1033 ( .A(n1196), .B(n474), .S(n604), .Z(n3065) );
  MUX2_X1 U1034 ( .A(n1197), .B(n477), .S(n603), .Z(n3064) );
  MUX2_X1 U1035 ( .A(n1198), .B(n480), .S(n603), .Z(n3063) );
  MUX2_X1 U1036 ( .A(n1199), .B(n483), .S(n603), .Z(n3062) );
  MUX2_X1 U1037 ( .A(n1200), .B(n486), .S(n603), .Z(n3061) );
  MUX2_X1 U1038 ( .A(n1201), .B(n489), .S(n603), .Z(n3060) );
  MUX2_X1 U1039 ( .A(n1202), .B(n492), .S(n603), .Z(n3059) );
  MUX2_X1 U1040 ( .A(n1203), .B(n495), .S(n603), .Z(n3058) );
  MUX2_X1 U1041 ( .A(n1204), .B(n498), .S(n603), .Z(n3057) );
  MUX2_X1 U1042 ( .A(n1205), .B(n501), .S(n603), .Z(n3056) );
  MUX2_X1 U1043 ( .A(n1206), .B(n504), .S(n603), .Z(n3055) );
  MUX2_X1 U1044 ( .A(n1207), .B(n507), .S(n603), .Z(n3054) );
  MUX2_X1 U1045 ( .A(n1208), .B(n510), .S(n603), .Z(n3053) );
  MUX2_X1 U1046 ( .A(n1209), .B(n513), .S(n602), .Z(n3052) );
  MUX2_X1 U1047 ( .A(n1210), .B(n516), .S(n602), .Z(n3051) );
  MUX2_X1 U1048 ( .A(n1211), .B(n519), .S(n602), .Z(n3050) );
  MUX2_X1 U1049 ( .A(n1212), .B(n522), .S(n602), .Z(n3049) );
  MUX2_X1 U1050 ( .A(n1213), .B(n525), .S(n602), .Z(n3048) );
  MUX2_X1 U1051 ( .A(n1214), .B(n528), .S(n602), .Z(n3047) );
  MUX2_X1 U1052 ( .A(n1215), .B(n531), .S(n602), .Z(n3046) );
  MUX2_X1 U1053 ( .A(n1216), .B(n534), .S(n602), .Z(n3045) );
  MUX2_X1 U1054 ( .A(n1217), .B(n537), .S(n602), .Z(n3044) );
  MUX2_X1 U1055 ( .A(n1218), .B(n540), .S(n602), .Z(n3043) );
  MUX2_X1 U1056 ( .A(n1219), .B(n543), .S(n602), .Z(n3042) );
  MUX2_X1 U1057 ( .A(n1220), .B(n546), .S(n602), .Z(n3041) );
  OAI21_X1 U1058 ( .B1(n940), .B2(n1153), .A(RESET), .ZN(n1189) );
  NAND3_X1 U1059 ( .A1(n941), .A2(n942), .A3(n1221), .ZN(n1153) );
  MUX2_X1 U1060 ( .A(n3856), .B(n450), .S(n607), .Z(n3040) );
  MUX2_X1 U1061 ( .A(n3874), .B(n456), .S(n607), .Z(n3039) );
  MUX2_X1 U1062 ( .A(n3910), .B(n459), .S(n607), .Z(n3038) );
  MUX2_X1 U1063 ( .A(n3928), .B(n462), .S(n607), .Z(n3037) );
  MUX2_X1 U1064 ( .A(n3946), .B(n465), .S(n607), .Z(n3036) );
  MUX2_X1 U1065 ( .A(n3964), .B(n468), .S(n607), .Z(n3035) );
  MUX2_X1 U1066 ( .A(n3982), .B(n471), .S(n607), .Z(n3034) );
  MUX2_X1 U1067 ( .A(n4000), .B(n474), .S(n607), .Z(n3033) );
  MUX2_X1 U1068 ( .A(n4018), .B(n477), .S(n606), .Z(n3032) );
  MUX2_X1 U1069 ( .A(n4036), .B(n480), .S(n606), .Z(n3031) );
  MUX2_X1 U1070 ( .A(n4054), .B(n483), .S(n606), .Z(n3030) );
  MUX2_X1 U1071 ( .A(n4072), .B(n486), .S(n606), .Z(n3029) );
  MUX2_X1 U1072 ( .A(n4108), .B(n489), .S(n606), .Z(n3028) );
  MUX2_X1 U1073 ( .A(n4126), .B(n492), .S(n606), .Z(n3027) );
  MUX2_X1 U1074 ( .A(n4144), .B(n495), .S(n606), .Z(n3026) );
  MUX2_X1 U1075 ( .A(n4162), .B(n498), .S(n606), .Z(n3025) );
  MUX2_X1 U1076 ( .A(n4180), .B(n501), .S(n606), .Z(n3024) );
  MUX2_X1 U1077 ( .A(n4198), .B(n504), .S(n606), .Z(n3023) );
  MUX2_X1 U1078 ( .A(n4216), .B(n507), .S(n606), .Z(n3022) );
  MUX2_X1 U1079 ( .A(n4234), .B(n510), .S(n606), .Z(n3021) );
  MUX2_X1 U1080 ( .A(n4252), .B(n513), .S(n605), .Z(n3020) );
  MUX2_X1 U1081 ( .A(n4270), .B(n516), .S(n605), .Z(n3019) );
  MUX2_X1 U1082 ( .A(n3730), .B(n519), .S(n605), .Z(n3018) );
  MUX2_X1 U1083 ( .A(n3748), .B(n522), .S(n605), .Z(n3017) );
  MUX2_X1 U1084 ( .A(n3766), .B(n525), .S(n605), .Z(n3016) );
  MUX2_X1 U1085 ( .A(n3784), .B(n528), .S(n605), .Z(n3015) );
  MUX2_X1 U1086 ( .A(n3802), .B(n531), .S(n605), .Z(n3014) );
  MUX2_X1 U1087 ( .A(n3820), .B(n534), .S(n605), .Z(n3013) );
  MUX2_X1 U1088 ( .A(n3838), .B(n537), .S(n605), .Z(n3012) );
  MUX2_X1 U1089 ( .A(n3892), .B(n540), .S(n605), .Z(n3011) );
  MUX2_X1 U1090 ( .A(n4090), .B(n543), .S(n605), .Z(n3010) );
  MUX2_X1 U1091 ( .A(n4288), .B(n546), .S(n605), .Z(n3009) );
  OAI21_X1 U1092 ( .B1(n870), .B2(n1223), .A(n833), .ZN(n1222) );
  MUX2_X1 U1093 ( .A(n3857), .B(n450), .S(n610), .Z(n3008) );
  MUX2_X1 U1094 ( .A(n3875), .B(n456), .S(n610), .Z(n3007) );
  MUX2_X1 U1095 ( .A(n3911), .B(n459), .S(n610), .Z(n3006) );
  MUX2_X1 U1096 ( .A(n3929), .B(n462), .S(n610), .Z(n3005) );
  MUX2_X1 U1097 ( .A(n3947), .B(n465), .S(n610), .Z(n3004) );
  MUX2_X1 U1098 ( .A(n3965), .B(n468), .S(n610), .Z(n3003) );
  MUX2_X1 U1099 ( .A(n3983), .B(n471), .S(n610), .Z(n3002) );
  MUX2_X1 U1100 ( .A(n4001), .B(n474), .S(n610), .Z(n3001) );
  MUX2_X1 U1101 ( .A(n4019), .B(n477), .S(n609), .Z(n3000) );
  MUX2_X1 U1102 ( .A(n4037), .B(n480), .S(n609), .Z(n2999) );
  MUX2_X1 U1103 ( .A(n4055), .B(n483), .S(n609), .Z(n2998) );
  MUX2_X1 U1104 ( .A(n4073), .B(n486), .S(n609), .Z(n2997) );
  MUX2_X1 U1105 ( .A(n4109), .B(n489), .S(n609), .Z(n2996) );
  MUX2_X1 U1106 ( .A(n4127), .B(n492), .S(n609), .Z(n2995) );
  MUX2_X1 U1107 ( .A(n4145), .B(n495), .S(n609), .Z(n2994) );
  MUX2_X1 U1108 ( .A(n4163), .B(n498), .S(n609), .Z(n2993) );
  MUX2_X1 U1109 ( .A(n4181), .B(n501), .S(n609), .Z(n2992) );
  MUX2_X1 U1110 ( .A(n4199), .B(n504), .S(n609), .Z(n2991) );
  MUX2_X1 U1111 ( .A(n4217), .B(n507), .S(n609), .Z(n2990) );
  MUX2_X1 U1112 ( .A(n4235), .B(n510), .S(n609), .Z(n2989) );
  MUX2_X1 U1113 ( .A(n4253), .B(n513), .S(n608), .Z(n2988) );
  MUX2_X1 U1114 ( .A(n4271), .B(n516), .S(n608), .Z(n2987) );
  MUX2_X1 U1115 ( .A(n3731), .B(n519), .S(n608), .Z(n2986) );
  MUX2_X1 U1116 ( .A(n3749), .B(n522), .S(n608), .Z(n2985) );
  MUX2_X1 U1117 ( .A(n3767), .B(n525), .S(n608), .Z(n2984) );
  MUX2_X1 U1118 ( .A(n3785), .B(n528), .S(n608), .Z(n2983) );
  MUX2_X1 U1119 ( .A(n3803), .B(n531), .S(n608), .Z(n2982) );
  MUX2_X1 U1120 ( .A(n3821), .B(n534), .S(n608), .Z(n2981) );
  MUX2_X1 U1121 ( .A(n3839), .B(n537), .S(n608), .Z(n2980) );
  MUX2_X1 U1122 ( .A(n3893), .B(n540), .S(n608), .Z(n2979) );
  MUX2_X1 U1123 ( .A(n4091), .B(n543), .S(n608), .Z(n2978) );
  MUX2_X1 U1124 ( .A(n4289), .B(n546), .S(n608), .Z(n2977) );
  OAI21_X1 U1125 ( .B1(n872), .B2(n1223), .A(RESET), .ZN(n1224) );
  MUX2_X1 U1126 ( .A(n1225), .B(n451), .S(n613), .Z(n2976) );
  MUX2_X1 U1127 ( .A(n1227), .B(n457), .S(n613), .Z(n2975) );
  MUX2_X1 U1128 ( .A(n1228), .B(n460), .S(n613), .Z(n2974) );
  MUX2_X1 U1129 ( .A(n1229), .B(n463), .S(n613), .Z(n2973) );
  MUX2_X1 U1130 ( .A(n1230), .B(n466), .S(n613), .Z(n2972) );
  MUX2_X1 U1131 ( .A(n1231), .B(n469), .S(n613), .Z(n2971) );
  MUX2_X1 U1132 ( .A(n1232), .B(n472), .S(n613), .Z(n2970) );
  MUX2_X1 U1133 ( .A(n1233), .B(n475), .S(n613), .Z(n2969) );
  MUX2_X1 U1134 ( .A(n1234), .B(n478), .S(n612), .Z(n2968) );
  MUX2_X1 U1135 ( .A(n1235), .B(n481), .S(n612), .Z(n2967) );
  MUX2_X1 U1136 ( .A(n1236), .B(n484), .S(n612), .Z(n2966) );
  MUX2_X1 U1137 ( .A(n1237), .B(n487), .S(n612), .Z(n2965) );
  MUX2_X1 U1138 ( .A(n1238), .B(n490), .S(n612), .Z(n2964) );
  MUX2_X1 U1139 ( .A(n1239), .B(n493), .S(n612), .Z(n2963) );
  MUX2_X1 U1140 ( .A(n1240), .B(n496), .S(n612), .Z(n2962) );
  MUX2_X1 U1141 ( .A(n1241), .B(n499), .S(n612), .Z(n2961) );
  MUX2_X1 U1142 ( .A(n1242), .B(n502), .S(n612), .Z(n2960) );
  MUX2_X1 U1143 ( .A(n1243), .B(n505), .S(n612), .Z(n2959) );
  MUX2_X1 U1144 ( .A(n1244), .B(n508), .S(n612), .Z(n2958) );
  MUX2_X1 U1145 ( .A(n1245), .B(n511), .S(n612), .Z(n2957) );
  MUX2_X1 U1146 ( .A(n1246), .B(n514), .S(n611), .Z(n2956) );
  MUX2_X1 U1147 ( .A(n1247), .B(n517), .S(n611), .Z(n2955) );
  MUX2_X1 U1148 ( .A(n1248), .B(n520), .S(n611), .Z(n2954) );
  MUX2_X1 U1149 ( .A(n1249), .B(n523), .S(n611), .Z(n2953) );
  MUX2_X1 U1150 ( .A(n1250), .B(n526), .S(n611), .Z(n2952) );
  MUX2_X1 U1151 ( .A(n1251), .B(n529), .S(n611), .Z(n2951) );
  MUX2_X1 U1152 ( .A(n1252), .B(n532), .S(n611), .Z(n2950) );
  MUX2_X1 U1153 ( .A(n1253), .B(n535), .S(n611), .Z(n2949) );
  MUX2_X1 U1154 ( .A(n1254), .B(n538), .S(n611), .Z(n2948) );
  MUX2_X1 U1155 ( .A(n1255), .B(n541), .S(n611), .Z(n2947) );
  MUX2_X1 U1156 ( .A(n1256), .B(n544), .S(n611), .Z(n2946) );
  MUX2_X1 U1157 ( .A(n1257), .B(n547), .S(n611), .Z(n2945) );
  OAI21_X1 U1158 ( .B1(n906), .B2(n1223), .A(n833), .ZN(n1226) );
  MUX2_X1 U1159 ( .A(n1258), .B(n451), .S(n616), .Z(n2944) );
  MUX2_X1 U1160 ( .A(n1260), .B(n457), .S(n616), .Z(n2943) );
  MUX2_X1 U1161 ( .A(n1261), .B(n460), .S(n616), .Z(n2942) );
  MUX2_X1 U1162 ( .A(n1262), .B(n463), .S(n616), .Z(n2941) );
  MUX2_X1 U1163 ( .A(n1263), .B(n466), .S(n616), .Z(n2940) );
  MUX2_X1 U1164 ( .A(n1264), .B(n469), .S(n616), .Z(n2939) );
  MUX2_X1 U1165 ( .A(n1265), .B(n472), .S(n616), .Z(n2938) );
  MUX2_X1 U1166 ( .A(n1266), .B(n475), .S(n616), .Z(n2937) );
  MUX2_X1 U1167 ( .A(n1267), .B(n478), .S(n615), .Z(n2936) );
  MUX2_X1 U1168 ( .A(n1268), .B(n481), .S(n615), .Z(n2935) );
  MUX2_X1 U1169 ( .A(n1269), .B(n484), .S(n615), .Z(n2934) );
  MUX2_X1 U1170 ( .A(n1270), .B(n487), .S(n615), .Z(n2933) );
  MUX2_X1 U1171 ( .A(n1271), .B(n490), .S(n615), .Z(n2932) );
  MUX2_X1 U1172 ( .A(n1272), .B(n493), .S(n615), .Z(n2931) );
  MUX2_X1 U1173 ( .A(n1273), .B(n496), .S(n615), .Z(n2930) );
  MUX2_X1 U1174 ( .A(n1274), .B(n499), .S(n615), .Z(n2929) );
  MUX2_X1 U1175 ( .A(n1275), .B(n502), .S(n615), .Z(n2928) );
  MUX2_X1 U1176 ( .A(n1276), .B(n505), .S(n615), .Z(n2927) );
  MUX2_X1 U1177 ( .A(n1277), .B(n508), .S(n615), .Z(n2926) );
  MUX2_X1 U1178 ( .A(n1278), .B(n511), .S(n615), .Z(n2925) );
  MUX2_X1 U1179 ( .A(n1279), .B(n514), .S(n614), .Z(n2924) );
  MUX2_X1 U1180 ( .A(n1280), .B(n517), .S(n614), .Z(n2923) );
  MUX2_X1 U1181 ( .A(n1281), .B(n520), .S(n614), .Z(n2922) );
  MUX2_X1 U1182 ( .A(n1282), .B(n523), .S(n614), .Z(n2921) );
  MUX2_X1 U1183 ( .A(n1283), .B(n526), .S(n614), .Z(n2920) );
  MUX2_X1 U1184 ( .A(n1284), .B(n529), .S(n614), .Z(n2919) );
  MUX2_X1 U1185 ( .A(n1285), .B(n532), .S(n614), .Z(n2918) );
  MUX2_X1 U1186 ( .A(n1286), .B(n535), .S(n614), .Z(n2917) );
  MUX2_X1 U1187 ( .A(n1287), .B(n538), .S(n614), .Z(n2916) );
  MUX2_X1 U1188 ( .A(n1288), .B(n541), .S(n614), .Z(n2915) );
  MUX2_X1 U1189 ( .A(n1289), .B(n544), .S(n614), .Z(n2914) );
  MUX2_X1 U1190 ( .A(n1290), .B(n547), .S(n614), .Z(n2913) );
  OAI21_X1 U1191 ( .B1(n940), .B2(n1223), .A(RESET), .ZN(n1259) );
  NAND3_X1 U1192 ( .A1(ADD_WR[2]), .A2(n942), .A3(n1221), .ZN(n1223) );
  INV_X1 U1193 ( .A(ADD_WR[3]), .ZN(n942) );
  MUX2_X1 U1194 ( .A(n3861), .B(n451), .S(n619), .Z(n2912) );
  MUX2_X1 U1195 ( .A(n3879), .B(n457), .S(n619), .Z(n2911) );
  MUX2_X1 U1196 ( .A(n3915), .B(n460), .S(n619), .Z(n2910) );
  MUX2_X1 U1197 ( .A(n3933), .B(n463), .S(n619), .Z(n2909) );
  MUX2_X1 U1198 ( .A(n3951), .B(n466), .S(n619), .Z(n2908) );
  MUX2_X1 U1199 ( .A(n3969), .B(n469), .S(n619), .Z(n2907) );
  MUX2_X1 U1200 ( .A(n3987), .B(n472), .S(n619), .Z(n2906) );
  MUX2_X1 U1201 ( .A(n4005), .B(n475), .S(n619), .Z(n2905) );
  MUX2_X1 U1202 ( .A(n4023), .B(n478), .S(n618), .Z(n2904) );
  MUX2_X1 U1203 ( .A(n4041), .B(n481), .S(n618), .Z(n2903) );
  MUX2_X1 U1204 ( .A(n4059), .B(n484), .S(n618), .Z(n2902) );
  MUX2_X1 U1205 ( .A(n4077), .B(n487), .S(n618), .Z(n2901) );
  MUX2_X1 U1206 ( .A(n4113), .B(n490), .S(n618), .Z(n2900) );
  MUX2_X1 U1207 ( .A(n4131), .B(n493), .S(n618), .Z(n2899) );
  MUX2_X1 U1208 ( .A(n4149), .B(n496), .S(n618), .Z(n2898) );
  MUX2_X1 U1209 ( .A(n4167), .B(n499), .S(n618), .Z(n2897) );
  MUX2_X1 U1210 ( .A(n4185), .B(n502), .S(n618), .Z(n2896) );
  MUX2_X1 U1211 ( .A(n4203), .B(n505), .S(n618), .Z(n2895) );
  MUX2_X1 U1212 ( .A(n4221), .B(n508), .S(n618), .Z(n2894) );
  MUX2_X1 U1213 ( .A(n4239), .B(n511), .S(n618), .Z(n2893) );
  MUX2_X1 U1214 ( .A(n4257), .B(n514), .S(n617), .Z(n2892) );
  MUX2_X1 U1215 ( .A(n4275), .B(n517), .S(n617), .Z(n2891) );
  MUX2_X1 U1216 ( .A(n3735), .B(n520), .S(n617), .Z(n2890) );
  MUX2_X1 U1217 ( .A(n3753), .B(n523), .S(n617), .Z(n2889) );
  MUX2_X1 U1218 ( .A(n3771), .B(n526), .S(n617), .Z(n2888) );
  MUX2_X1 U1219 ( .A(n3789), .B(n529), .S(n617), .Z(n2887) );
  MUX2_X1 U1220 ( .A(n3807), .B(n532), .S(n617), .Z(n2886) );
  MUX2_X1 U1221 ( .A(n3825), .B(n535), .S(n617), .Z(n2885) );
  MUX2_X1 U1222 ( .A(n3843), .B(n538), .S(n617), .Z(n2884) );
  MUX2_X1 U1223 ( .A(n3897), .B(n541), .S(n617), .Z(n2883) );
  MUX2_X1 U1224 ( .A(n4095), .B(n544), .S(n617), .Z(n2882) );
  MUX2_X1 U1225 ( .A(n4293), .B(n547), .S(n617), .Z(n2881) );
  OAI21_X1 U1226 ( .B1(n870), .B2(n1292), .A(RESET), .ZN(n1291) );
  MUX2_X1 U1227 ( .A(n3860), .B(n451), .S(n622), .Z(n2880) );
  MUX2_X1 U1228 ( .A(n3878), .B(n457), .S(n622), .Z(n2879) );
  MUX2_X1 U1229 ( .A(n3914), .B(n460), .S(n622), .Z(n2878) );
  MUX2_X1 U1230 ( .A(n3932), .B(n463), .S(n622), .Z(n2877) );
  MUX2_X1 U1231 ( .A(n3950), .B(n466), .S(n622), .Z(n2876) );
  MUX2_X1 U1232 ( .A(n3968), .B(n469), .S(n622), .Z(n2875) );
  MUX2_X1 U1233 ( .A(n3986), .B(n472), .S(n622), .Z(n2874) );
  MUX2_X1 U1234 ( .A(n4004), .B(n475), .S(n622), .Z(n2873) );
  MUX2_X1 U1235 ( .A(n4022), .B(n478), .S(n621), .Z(n2872) );
  MUX2_X1 U1236 ( .A(n4040), .B(n481), .S(n621), .Z(n2871) );
  MUX2_X1 U1237 ( .A(n4058), .B(n484), .S(n621), .Z(n2870) );
  MUX2_X1 U1238 ( .A(n4076), .B(n487), .S(n621), .Z(n2869) );
  MUX2_X1 U1239 ( .A(n4112), .B(n490), .S(n621), .Z(n2868) );
  MUX2_X1 U1240 ( .A(n4130), .B(n493), .S(n621), .Z(n2867) );
  MUX2_X1 U1241 ( .A(n4148), .B(n496), .S(n621), .Z(n2866) );
  MUX2_X1 U1242 ( .A(n4166), .B(n499), .S(n621), .Z(n2865) );
  MUX2_X1 U1243 ( .A(n4184), .B(n502), .S(n621), .Z(n2864) );
  MUX2_X1 U1244 ( .A(n4202), .B(n505), .S(n621), .Z(n2863) );
  MUX2_X1 U1245 ( .A(n4220), .B(n508), .S(n621), .Z(n2862) );
  MUX2_X1 U1246 ( .A(n4238), .B(n511), .S(n621), .Z(n2861) );
  MUX2_X1 U1247 ( .A(n4256), .B(n514), .S(n620), .Z(n2860) );
  MUX2_X1 U1248 ( .A(n4274), .B(n517), .S(n620), .Z(n2859) );
  MUX2_X1 U1249 ( .A(n3734), .B(n520), .S(n620), .Z(n2858) );
  MUX2_X1 U1250 ( .A(n3752), .B(n523), .S(n620), .Z(n2857) );
  MUX2_X1 U1251 ( .A(n3770), .B(n526), .S(n620), .Z(n2856) );
  MUX2_X1 U1252 ( .A(n3788), .B(n529), .S(n620), .Z(n2855) );
  MUX2_X1 U1253 ( .A(n3806), .B(n532), .S(n620), .Z(n2854) );
  MUX2_X1 U1254 ( .A(n3824), .B(n535), .S(n620), .Z(n2853) );
  MUX2_X1 U1255 ( .A(n3842), .B(n538), .S(n620), .Z(n2852) );
  MUX2_X1 U1256 ( .A(n3896), .B(n541), .S(n620), .Z(n2851) );
  MUX2_X1 U1257 ( .A(n4094), .B(n544), .S(n620), .Z(n2850) );
  MUX2_X1 U1258 ( .A(n4292), .B(n547), .S(n620), .Z(n2849) );
  OAI21_X1 U1259 ( .B1(n872), .B2(n1292), .A(RESET), .ZN(n1293) );
  MUX2_X1 U1260 ( .A(n1294), .B(n451), .S(n625), .Z(n2848) );
  MUX2_X1 U1261 ( .A(n1296), .B(n457), .S(n625), .Z(n2847) );
  MUX2_X1 U1262 ( .A(n1297), .B(n460), .S(n625), .Z(n2846) );
  MUX2_X1 U1263 ( .A(n1298), .B(n463), .S(n625), .Z(n2845) );
  MUX2_X1 U1264 ( .A(n1299), .B(n466), .S(n625), .Z(n2844) );
  MUX2_X1 U1265 ( .A(n1300), .B(n469), .S(n625), .Z(n2843) );
  MUX2_X1 U1266 ( .A(n1301), .B(n472), .S(n625), .Z(n2842) );
  MUX2_X1 U1267 ( .A(n1302), .B(n475), .S(n625), .Z(n2841) );
  MUX2_X1 U1268 ( .A(n1303), .B(n478), .S(n624), .Z(n2840) );
  MUX2_X1 U1269 ( .A(n1304), .B(n481), .S(n624), .Z(n2839) );
  MUX2_X1 U1270 ( .A(n1305), .B(n484), .S(n624), .Z(n2838) );
  MUX2_X1 U1271 ( .A(n1306), .B(n487), .S(n624), .Z(n2837) );
  MUX2_X1 U1272 ( .A(n1307), .B(n490), .S(n624), .Z(n2836) );
  MUX2_X1 U1273 ( .A(n1308), .B(n493), .S(n624), .Z(n2835) );
  MUX2_X1 U1274 ( .A(n1309), .B(n496), .S(n624), .Z(n2834) );
  MUX2_X1 U1275 ( .A(n1310), .B(n499), .S(n624), .Z(n2833) );
  MUX2_X1 U1276 ( .A(n1311), .B(n502), .S(n624), .Z(n2832) );
  MUX2_X1 U1277 ( .A(n1312), .B(n505), .S(n624), .Z(n2831) );
  MUX2_X1 U1278 ( .A(n1313), .B(n508), .S(n624), .Z(n2830) );
  MUX2_X1 U1279 ( .A(n1314), .B(n511), .S(n624), .Z(n2829) );
  MUX2_X1 U1280 ( .A(n1315), .B(n514), .S(n623), .Z(n2828) );
  MUX2_X1 U1281 ( .A(n1316), .B(n517), .S(n623), .Z(n2827) );
  MUX2_X1 U1282 ( .A(n1317), .B(n520), .S(n623), .Z(n2826) );
  MUX2_X1 U1283 ( .A(n1318), .B(n523), .S(n623), .Z(n2825) );
  MUX2_X1 U1284 ( .A(n1319), .B(n526), .S(n623), .Z(n2824) );
  MUX2_X1 U1285 ( .A(n1320), .B(n529), .S(n623), .Z(n2823) );
  MUX2_X1 U1286 ( .A(n1321), .B(n532), .S(n623), .Z(n2822) );
  MUX2_X1 U1287 ( .A(n1322), .B(n535), .S(n623), .Z(n2821) );
  MUX2_X1 U1288 ( .A(n1323), .B(n538), .S(n623), .Z(n2820) );
  MUX2_X1 U1289 ( .A(n1324), .B(n541), .S(n623), .Z(n2819) );
  MUX2_X1 U1290 ( .A(n1325), .B(n544), .S(n623), .Z(n2818) );
  MUX2_X1 U1291 ( .A(n1326), .B(n547), .S(n623), .Z(n2817) );
  OAI21_X1 U1292 ( .B1(n906), .B2(n1292), .A(RESET), .ZN(n1295) );
  MUX2_X1 U1293 ( .A(n1327), .B(n451), .S(n628), .Z(n2816) );
  MUX2_X1 U1294 ( .A(n1329), .B(n457), .S(n628), .Z(n2815) );
  MUX2_X1 U1295 ( .A(n1330), .B(n460), .S(n628), .Z(n2814) );
  MUX2_X1 U1296 ( .A(n1331), .B(n463), .S(n628), .Z(n2813) );
  MUX2_X1 U1297 ( .A(n1332), .B(n466), .S(n628), .Z(n2812) );
  MUX2_X1 U1298 ( .A(n1333), .B(n469), .S(n628), .Z(n2811) );
  MUX2_X1 U1299 ( .A(n1334), .B(n472), .S(n628), .Z(n2810) );
  MUX2_X1 U1300 ( .A(n1335), .B(n475), .S(n628), .Z(n2809) );
  MUX2_X1 U1301 ( .A(n1336), .B(n478), .S(n627), .Z(n2808) );
  MUX2_X1 U1302 ( .A(n1337), .B(n481), .S(n627), .Z(n2807) );
  MUX2_X1 U1303 ( .A(n1338), .B(n484), .S(n627), .Z(n2806) );
  MUX2_X1 U1304 ( .A(n1339), .B(n487), .S(n627), .Z(n2805) );
  MUX2_X1 U1305 ( .A(n1340), .B(n490), .S(n627), .Z(n2804) );
  MUX2_X1 U1306 ( .A(n1341), .B(n493), .S(n627), .Z(n2803) );
  MUX2_X1 U1307 ( .A(n1342), .B(n496), .S(n627), .Z(n2802) );
  MUX2_X1 U1308 ( .A(n1343), .B(n499), .S(n627), .Z(n2801) );
  MUX2_X1 U1309 ( .A(n1344), .B(n502), .S(n627), .Z(n2800) );
  MUX2_X1 U1310 ( .A(n1345), .B(n505), .S(n627), .Z(n2799) );
  MUX2_X1 U1311 ( .A(n1346), .B(n508), .S(n627), .Z(n2798) );
  MUX2_X1 U1312 ( .A(n1347), .B(n511), .S(n627), .Z(n2797) );
  MUX2_X1 U1313 ( .A(n1348), .B(n514), .S(n626), .Z(n2796) );
  MUX2_X1 U1314 ( .A(n1349), .B(n517), .S(n626), .Z(n2795) );
  MUX2_X1 U1315 ( .A(n1350), .B(n520), .S(n626), .Z(n2794) );
  MUX2_X1 U1316 ( .A(n1351), .B(n523), .S(n626), .Z(n2793) );
  MUX2_X1 U1317 ( .A(n1352), .B(n526), .S(n626), .Z(n2792) );
  MUX2_X1 U1318 ( .A(n1353), .B(n529), .S(n626), .Z(n2791) );
  MUX2_X1 U1319 ( .A(n1354), .B(n532), .S(n626), .Z(n2790) );
  MUX2_X1 U1320 ( .A(n1355), .B(n535), .S(n626), .Z(n2789) );
  MUX2_X1 U1321 ( .A(n1356), .B(n538), .S(n626), .Z(n2788) );
  MUX2_X1 U1322 ( .A(n1357), .B(n541), .S(n626), .Z(n2787) );
  MUX2_X1 U1323 ( .A(n1358), .B(n544), .S(n626), .Z(n2786) );
  MUX2_X1 U1324 ( .A(n1359), .B(n547), .S(n626), .Z(n2785) );
  OAI21_X1 U1325 ( .B1(n940), .B2(n1292), .A(RESET), .ZN(n1328) );
  NAND3_X1 U1326 ( .A1(ADD_WR[3]), .A2(n941), .A3(n1221), .ZN(n1292) );
  INV_X1 U1327 ( .A(ADD_WR[2]), .ZN(n941) );
  MUX2_X1 U1328 ( .A(n1360), .B(n451), .S(n631), .Z(n2784) );
  MUX2_X1 U1329 ( .A(n1362), .B(n457), .S(n631), .Z(n2783) );
  MUX2_X1 U1330 ( .A(n1363), .B(n460), .S(n631), .Z(n2782) );
  MUX2_X1 U1331 ( .A(n1364), .B(n463), .S(n631), .Z(n2781) );
  MUX2_X1 U1332 ( .A(n1365), .B(n466), .S(n631), .Z(n2780) );
  MUX2_X1 U1333 ( .A(n1366), .B(n469), .S(n631), .Z(n2779) );
  MUX2_X1 U1334 ( .A(n1367), .B(n472), .S(n631), .Z(n2778) );
  MUX2_X1 U1335 ( .A(n1368), .B(n475), .S(n631), .Z(n2777) );
  MUX2_X1 U1336 ( .A(n1369), .B(n478), .S(n630), .Z(n2776) );
  MUX2_X1 U1337 ( .A(n1370), .B(n481), .S(n630), .Z(n2775) );
  MUX2_X1 U1338 ( .A(n1371), .B(n484), .S(n630), .Z(n2774) );
  MUX2_X1 U1339 ( .A(n1372), .B(n487), .S(n630), .Z(n2773) );
  MUX2_X1 U1340 ( .A(n1373), .B(n490), .S(n630), .Z(n2772) );
  MUX2_X1 U1341 ( .A(n1374), .B(n493), .S(n630), .Z(n2771) );
  MUX2_X1 U1342 ( .A(n1375), .B(n496), .S(n630), .Z(n2770) );
  MUX2_X1 U1343 ( .A(n1376), .B(n499), .S(n630), .Z(n2769) );
  MUX2_X1 U1344 ( .A(n1377), .B(n502), .S(n630), .Z(n2768) );
  MUX2_X1 U1345 ( .A(n1378), .B(n505), .S(n630), .Z(n2767) );
  MUX2_X1 U1346 ( .A(n1379), .B(n508), .S(n630), .Z(n2766) );
  MUX2_X1 U1347 ( .A(n1380), .B(n511), .S(n630), .Z(n2765) );
  MUX2_X1 U1348 ( .A(n1381), .B(n514), .S(n629), .Z(n2764) );
  MUX2_X1 U1349 ( .A(n1382), .B(n517), .S(n629), .Z(n2763) );
  MUX2_X1 U1350 ( .A(n1383), .B(n520), .S(n629), .Z(n2762) );
  MUX2_X1 U1351 ( .A(n1384), .B(n523), .S(n629), .Z(n2761) );
  MUX2_X1 U1352 ( .A(n1385), .B(n526), .S(n629), .Z(n2760) );
  MUX2_X1 U1353 ( .A(n1386), .B(n529), .S(n629), .Z(n2759) );
  MUX2_X1 U1354 ( .A(n1387), .B(n532), .S(n629), .Z(n2758) );
  MUX2_X1 U1355 ( .A(n1388), .B(n535), .S(n629), .Z(n2757) );
  MUX2_X1 U1356 ( .A(n1389), .B(n538), .S(n629), .Z(n2756) );
  MUX2_X1 U1357 ( .A(n1390), .B(n541), .S(n629), .Z(n2755) );
  MUX2_X1 U1358 ( .A(n1391), .B(n544), .S(n629), .Z(n2754) );
  MUX2_X1 U1359 ( .A(n1392), .B(n547), .S(n629), .Z(n2753) );
  OAI21_X1 U1360 ( .B1(n870), .B2(n1393), .A(RESET), .ZN(n1361) );
  NAND2_X1 U1361 ( .A1(n1394), .A2(n1395), .ZN(n870) );
  MUX2_X1 U1362 ( .A(n1396), .B(n451), .S(n634), .Z(n2752) );
  MUX2_X1 U1363 ( .A(n1398), .B(n457), .S(n634), .Z(n2751) );
  MUX2_X1 U1364 ( .A(n1399), .B(n460), .S(n634), .Z(n2750) );
  MUX2_X1 U1365 ( .A(n1400), .B(n463), .S(n634), .Z(n2749) );
  MUX2_X1 U1366 ( .A(n1401), .B(n466), .S(n634), .Z(n2748) );
  MUX2_X1 U1367 ( .A(n1402), .B(n469), .S(n634), .Z(n2747) );
  MUX2_X1 U1368 ( .A(n1403), .B(n472), .S(n634), .Z(n2746) );
  MUX2_X1 U1369 ( .A(n1404), .B(n475), .S(n634), .Z(n2745) );
  MUX2_X1 U1370 ( .A(n1405), .B(n478), .S(n633), .Z(n2744) );
  MUX2_X1 U1371 ( .A(n1406), .B(n481), .S(n633), .Z(n2743) );
  MUX2_X1 U1372 ( .A(n1407), .B(n484), .S(n633), .Z(n2742) );
  MUX2_X1 U1373 ( .A(n1408), .B(n487), .S(n633), .Z(n2741) );
  MUX2_X1 U1374 ( .A(n1409), .B(n490), .S(n633), .Z(n2740) );
  MUX2_X1 U1375 ( .A(n1410), .B(n493), .S(n633), .Z(n2739) );
  MUX2_X1 U1376 ( .A(n1411), .B(n496), .S(n633), .Z(n2738) );
  MUX2_X1 U1377 ( .A(n1412), .B(n499), .S(n633), .Z(n2737) );
  MUX2_X1 U1378 ( .A(n1413), .B(n502), .S(n633), .Z(n2736) );
  MUX2_X1 U1379 ( .A(n1414), .B(n505), .S(n633), .Z(n2735) );
  MUX2_X1 U1380 ( .A(n1415), .B(n508), .S(n633), .Z(n2734) );
  MUX2_X1 U1381 ( .A(n1416), .B(n511), .S(n633), .Z(n2733) );
  MUX2_X1 U1382 ( .A(n1417), .B(n514), .S(n632), .Z(n2732) );
  MUX2_X1 U1383 ( .A(n1418), .B(n517), .S(n632), .Z(n2731) );
  MUX2_X1 U1384 ( .A(n1419), .B(n520), .S(n632), .Z(n2730) );
  MUX2_X1 U1385 ( .A(n1420), .B(n523), .S(n632), .Z(n2729) );
  MUX2_X1 U1386 ( .A(n1421), .B(n526), .S(n632), .Z(n2728) );
  MUX2_X1 U1387 ( .A(n1422), .B(n529), .S(n632), .Z(n2727) );
  MUX2_X1 U1388 ( .A(n1423), .B(n532), .S(n632), .Z(n2726) );
  MUX2_X1 U1389 ( .A(n1424), .B(n535), .S(n632), .Z(n2725) );
  MUX2_X1 U1390 ( .A(n1425), .B(n538), .S(n632), .Z(n2724) );
  MUX2_X1 U1391 ( .A(n1426), .B(n541), .S(n632), .Z(n2723) );
  MUX2_X1 U1392 ( .A(n1427), .B(n544), .S(n632), .Z(n2722) );
  MUX2_X1 U1393 ( .A(n1428), .B(n547), .S(n632), .Z(n2721) );
  OAI21_X1 U1394 ( .B1(n872), .B2(n1393), .A(RESET), .ZN(n1397) );
  NAND2_X1 U1395 ( .A1(ADD_WR[0]), .A2(n1394), .ZN(n872) );
  INV_X1 U1396 ( .A(ADD_WR[1]), .ZN(n1394) );
  MUX2_X1 U1397 ( .A(n3865), .B(n451), .S(n637), .Z(n2720) );
  MUX2_X1 U1398 ( .A(n3883), .B(n457), .S(n637), .Z(n2719) );
  MUX2_X1 U1399 ( .A(n3919), .B(n460), .S(n637), .Z(n2718) );
  MUX2_X1 U1400 ( .A(n3937), .B(n463), .S(n637), .Z(n2717) );
  MUX2_X1 U1401 ( .A(n3955), .B(n466), .S(n637), .Z(n2716) );
  MUX2_X1 U1402 ( .A(n3973), .B(n469), .S(n637), .Z(n2715) );
  MUX2_X1 U1403 ( .A(n3991), .B(n472), .S(n637), .Z(n2714) );
  MUX2_X1 U1404 ( .A(n4009), .B(n475), .S(n637), .Z(n2713) );
  MUX2_X1 U1405 ( .A(n4027), .B(n478), .S(n636), .Z(n2712) );
  MUX2_X1 U1406 ( .A(n4045), .B(n481), .S(n636), .Z(n2711) );
  MUX2_X1 U1407 ( .A(n4063), .B(n484), .S(n636), .Z(n2710) );
  MUX2_X1 U1408 ( .A(n4081), .B(n487), .S(n636), .Z(n2709) );
  MUX2_X1 U1409 ( .A(n4117), .B(n490), .S(n636), .Z(n2708) );
  MUX2_X1 U1410 ( .A(n4135), .B(n493), .S(n636), .Z(n2707) );
  MUX2_X1 U1411 ( .A(n4153), .B(n496), .S(n636), .Z(n2706) );
  MUX2_X1 U1412 ( .A(n4171), .B(n499), .S(n636), .Z(n2705) );
  MUX2_X1 U1413 ( .A(n4189), .B(n502), .S(n636), .Z(n2704) );
  MUX2_X1 U1414 ( .A(n4207), .B(n505), .S(n636), .Z(n2703) );
  MUX2_X1 U1415 ( .A(n4225), .B(n508), .S(n636), .Z(n2702) );
  MUX2_X1 U1416 ( .A(n4243), .B(n511), .S(n636), .Z(n2701) );
  MUX2_X1 U1417 ( .A(n4261), .B(n514), .S(n635), .Z(n2700) );
  MUX2_X1 U1418 ( .A(n4279), .B(n517), .S(n635), .Z(n2699) );
  MUX2_X1 U1419 ( .A(n3739), .B(n520), .S(n635), .Z(n2698) );
  MUX2_X1 U1420 ( .A(n3757), .B(n523), .S(n635), .Z(n2697) );
  MUX2_X1 U1421 ( .A(n3775), .B(n526), .S(n635), .Z(n2696) );
  MUX2_X1 U1422 ( .A(n3793), .B(n529), .S(n635), .Z(n2695) );
  MUX2_X1 U1423 ( .A(n3811), .B(n532), .S(n635), .Z(n2694) );
  MUX2_X1 U1424 ( .A(n3829), .B(n535), .S(n635), .Z(n2693) );
  MUX2_X1 U1425 ( .A(n3847), .B(n538), .S(n635), .Z(n2692) );
  MUX2_X1 U1426 ( .A(n3901), .B(n541), .S(n635), .Z(n2691) );
  MUX2_X1 U1427 ( .A(n4099), .B(n544), .S(n635), .Z(n2690) );
  MUX2_X1 U1428 ( .A(n4297), .B(n547), .S(n635), .Z(n2689) );
  OAI21_X1 U1429 ( .B1(n906), .B2(n1393), .A(RESET), .ZN(n1429) );
  NAND2_X1 U1430 ( .A1(ADD_WR[1]), .A2(n1395), .ZN(n906) );
  INV_X1 U1431 ( .A(ADD_WR[0]), .ZN(n1395) );
  MUX2_X1 U1432 ( .A(n3864), .B(n451), .S(n640), .Z(n2688) );
  AND2_X1 U1433 ( .A1(RESET), .A2(DATAIN[31]), .ZN(n836) );
  MUX2_X1 U1434 ( .A(n3882), .B(n457), .S(n640), .Z(n2687) );
  AND2_X1 U1435 ( .A1(DATAIN[30]), .A2(RESET), .ZN(n838) );
  MUX2_X1 U1436 ( .A(n3918), .B(n460), .S(n640), .Z(n2686) );
  AND2_X1 U1437 ( .A1(DATAIN[29]), .A2(RESET), .ZN(n839) );
  MUX2_X1 U1438 ( .A(n3936), .B(n463), .S(n640), .Z(n2685) );
  AND2_X1 U1439 ( .A1(DATAIN[28]), .A2(n834), .ZN(n840) );
  MUX2_X1 U1440 ( .A(n3954), .B(n466), .S(n640), .Z(n2684) );
  AND2_X1 U1441 ( .A1(DATAIN[27]), .A2(n834), .ZN(n841) );
  MUX2_X1 U1442 ( .A(n3972), .B(n469), .S(n640), .Z(n2683) );
  AND2_X1 U1443 ( .A1(DATAIN[26]), .A2(n834), .ZN(n842) );
  MUX2_X1 U1444 ( .A(n3990), .B(n472), .S(n640), .Z(n2682) );
  AND2_X1 U1445 ( .A1(DATAIN[25]), .A2(RESET), .ZN(n843) );
  MUX2_X1 U1446 ( .A(n4008), .B(n475), .S(n640), .Z(n2681) );
  AND2_X1 U1447 ( .A1(DATAIN[24]), .A2(n834), .ZN(n844) );
  MUX2_X1 U1448 ( .A(n4026), .B(n478), .S(n639), .Z(n2680) );
  AND2_X1 U1449 ( .A1(DATAIN[23]), .A2(n834), .ZN(n845) );
  MUX2_X1 U1450 ( .A(n4044), .B(n481), .S(n639), .Z(n2679) );
  AND2_X1 U1451 ( .A1(DATAIN[22]), .A2(n834), .ZN(n846) );
  MUX2_X1 U1452 ( .A(n4062), .B(n484), .S(n639), .Z(n2678) );
  AND2_X1 U1453 ( .A1(DATAIN[21]), .A2(n834), .ZN(n847) );
  MUX2_X1 U1454 ( .A(n4080), .B(n487), .S(n639), .Z(n2677) );
  AND2_X1 U1455 ( .A1(DATAIN[20]), .A2(n834), .ZN(n848) );
  MUX2_X1 U1456 ( .A(n4116), .B(n490), .S(n639), .Z(n2676) );
  AND2_X1 U1457 ( .A1(DATAIN[19]), .A2(n834), .ZN(n849) );
  MUX2_X1 U1458 ( .A(n4134), .B(n493), .S(n639), .Z(n2675) );
  AND2_X1 U1459 ( .A1(DATAIN[18]), .A2(n834), .ZN(n850) );
  MUX2_X1 U1460 ( .A(n4152), .B(n496), .S(n639), .Z(n2674) );
  AND2_X1 U1461 ( .A1(DATAIN[17]), .A2(n834), .ZN(n851) );
  MUX2_X1 U1462 ( .A(n4170), .B(n499), .S(n639), .Z(n2673) );
  AND2_X1 U1463 ( .A1(DATAIN[16]), .A2(n834), .ZN(n852) );
  MUX2_X1 U1464 ( .A(n4188), .B(n502), .S(n639), .Z(n2672) );
  AND2_X1 U1465 ( .A1(DATAIN[15]), .A2(n834), .ZN(n853) );
  MUX2_X1 U1466 ( .A(n4206), .B(n505), .S(n639), .Z(n2671) );
  AND2_X1 U1467 ( .A1(DATAIN[14]), .A2(n834), .ZN(n854) );
  MUX2_X1 U1468 ( .A(n4224), .B(n508), .S(n639), .Z(n2670) );
  AND2_X1 U1469 ( .A1(DATAIN[13]), .A2(n834), .ZN(n855) );
  MUX2_X1 U1470 ( .A(n4242), .B(n511), .S(n639), .Z(n2669) );
  AND2_X1 U1471 ( .A1(DATAIN[12]), .A2(n834), .ZN(n856) );
  MUX2_X1 U1472 ( .A(n4260), .B(n514), .S(n638), .Z(n2668) );
  AND2_X1 U1473 ( .A1(DATAIN[11]), .A2(n834), .ZN(n857) );
  MUX2_X1 U1474 ( .A(n4278), .B(n517), .S(n638), .Z(n2667) );
  AND2_X1 U1475 ( .A1(DATAIN[10]), .A2(n834), .ZN(n858) );
  MUX2_X1 U1476 ( .A(n3738), .B(n520), .S(n638), .Z(n2666) );
  AND2_X1 U1477 ( .A1(DATAIN[9]), .A2(n834), .ZN(n859) );
  MUX2_X1 U1478 ( .A(n3756), .B(n523), .S(n638), .Z(n2665) );
  AND2_X1 U1479 ( .A1(DATAIN[8]), .A2(n834), .ZN(n860) );
  MUX2_X1 U1480 ( .A(n3774), .B(n526), .S(n638), .Z(n2664) );
  AND2_X1 U1481 ( .A1(DATAIN[7]), .A2(n834), .ZN(n861) );
  MUX2_X1 U1482 ( .A(n3792), .B(n529), .S(n638), .Z(n2663) );
  AND2_X1 U1483 ( .A1(DATAIN[6]), .A2(n834), .ZN(n862) );
  MUX2_X1 U1484 ( .A(n3810), .B(n532), .S(n638), .Z(n2662) );
  AND2_X1 U1485 ( .A1(DATAIN[5]), .A2(RESET), .ZN(n863) );
  MUX2_X1 U1486 ( .A(n3828), .B(n535), .S(n638), .Z(n2661) );
  AND2_X1 U1487 ( .A1(DATAIN[4]), .A2(RESET), .ZN(n864) );
  MUX2_X1 U1488 ( .A(n3846), .B(n538), .S(n638), .Z(n2660) );
  AND2_X1 U1489 ( .A1(DATAIN[3]), .A2(RESET), .ZN(n865) );
  MUX2_X1 U1490 ( .A(n3900), .B(n541), .S(n638), .Z(n2659) );
  AND2_X1 U1491 ( .A1(DATAIN[2]), .A2(RESET), .ZN(n866) );
  MUX2_X1 U1492 ( .A(n4098), .B(n544), .S(n638), .Z(n2658) );
  AND2_X1 U1493 ( .A1(DATAIN[1]), .A2(RESET), .ZN(n867) );
  MUX2_X1 U1494 ( .A(n4296), .B(n547), .S(n638), .Z(n2657) );
  OAI21_X1 U1495 ( .B1(n940), .B2(n1393), .A(RESET), .ZN(n1430) );
  NAND3_X1 U1496 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .A3(n1221), .ZN(n1393) );
  AND2_X1 U1497 ( .A1(ADD_WR[4]), .A2(WR), .ZN(n1221) );
  NAND2_X1 U1498 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .ZN(n940) );
  AND2_X1 U1499 ( .A1(DATAIN[0]), .A2(n834), .ZN(n868) );
  NAND2_X1 U1500 ( .A1(n1431), .A2(n1432), .ZN(OUT2[9]) );
  NOR4_X1 U1501 ( .A1(n1433), .A2(n1434), .A3(n1435), .A4(n1436), .ZN(n1432)
         );
  OAI221_X1 U1502 ( .B1(n1), .B2(n643), .C1(n225), .C2(n646), .A(n1439), .ZN(
        n1436) );
  AOI22_X1 U1503 ( .A1(n649), .A2(n930), .B1(n652), .B2(n896), .ZN(n1439) );
  OAI221_X1 U1504 ( .B1(n2), .B2(n655), .C1(n226), .C2(n658), .A(n1444), .ZN(
        n1435) );
  AOI22_X1 U1505 ( .A1(n661), .A2(n1003), .B1(n664), .B2(n970), .ZN(n1444) );
  OAI221_X1 U1506 ( .B1(n3), .B2(n667), .C1(n227), .C2(n670), .A(n1449), .ZN(
        n1434) );
  AOI22_X1 U1507 ( .A1(n673), .A2(n1072), .B1(n676), .B2(n1039), .ZN(n1449) );
  OAI221_X1 U1508 ( .B1(n4), .B2(n679), .C1(n228), .C2(n682), .A(n1454), .ZN(
        n1433) );
  AOI22_X1 U1509 ( .A1(n685), .A2(n1141), .B1(n688), .B2(n1108), .ZN(n1454) );
  NOR4_X1 U1510 ( .A1(n1457), .A2(n1458), .A3(n1459), .A4(n1460), .ZN(n1431)
         );
  OAI221_X1 U1511 ( .B1(n3736), .B2(n691), .C1(n3737), .C2(n694), .A(n1463), 
        .ZN(n1460) );
  AOI22_X1 U1512 ( .A1(n697), .A2(n3738), .B1(n700), .B2(n3739), .ZN(n1463) );
  OAI221_X1 U1513 ( .B1(n5), .B2(n703), .C1(n229), .C2(n706), .A(n1468), .ZN(
        n1459) );
  AOI22_X1 U1514 ( .A1(n709), .A2(n1317), .B1(n712), .B2(n1350), .ZN(n1468) );
  OAI221_X1 U1515 ( .B1(n6), .B2(n715), .C1(n230), .C2(n718), .A(n1473), .ZN(
        n1458) );
  AOI22_X1 U1516 ( .A1(n721), .A2(n1178), .B1(n724), .B2(n1211), .ZN(n1473) );
  OAI221_X1 U1517 ( .B1(n7), .B2(n727), .C1(n231), .C2(n730), .A(n1478), .ZN(
        n1457) );
  AOI22_X1 U1518 ( .A1(n733), .A2(n1248), .B1(n736), .B2(n1281), .ZN(n1478) );
  NAND2_X1 U1519 ( .A1(n1481), .A2(n1482), .ZN(OUT2[8]) );
  NOR4_X1 U1520 ( .A1(n1483), .A2(n1484), .A3(n1485), .A4(n1486), .ZN(n1482)
         );
  OAI221_X1 U1521 ( .B1(n8), .B2(n643), .C1(n232), .C2(n646), .A(n1487), .ZN(
        n1486) );
  AOI22_X1 U1522 ( .A1(n649), .A2(n931), .B1(n652), .B2(n897), .ZN(n1487) );
  OAI221_X1 U1523 ( .B1(n9), .B2(n655), .C1(n233), .C2(n658), .A(n1488), .ZN(
        n1485) );
  AOI22_X1 U1524 ( .A1(n661), .A2(n1004), .B1(n664), .B2(n971), .ZN(n1488) );
  OAI221_X1 U1525 ( .B1(n10), .B2(n667), .C1(n234), .C2(n670), .A(n1489), .ZN(
        n1484) );
  AOI22_X1 U1526 ( .A1(n673), .A2(n1073), .B1(n676), .B2(n1040), .ZN(n1489) );
  OAI221_X1 U1527 ( .B1(n11), .B2(n679), .C1(n235), .C2(n682), .A(n1490), .ZN(
        n1483) );
  AOI22_X1 U1528 ( .A1(n685), .A2(n1142), .B1(n688), .B2(n1109), .ZN(n1490) );
  NOR4_X1 U1529 ( .A1(n1491), .A2(n1492), .A3(n1493), .A4(n1494), .ZN(n1481)
         );
  OAI221_X1 U1530 ( .B1(n3754), .B2(n691), .C1(n3755), .C2(n694), .A(n1495), 
        .ZN(n1494) );
  AOI22_X1 U1531 ( .A1(n697), .A2(n3756), .B1(n700), .B2(n3757), .ZN(n1495) );
  OAI221_X1 U1532 ( .B1(n12), .B2(n703), .C1(n236), .C2(n706), .A(n1496), .ZN(
        n1493) );
  AOI22_X1 U1533 ( .A1(n709), .A2(n1318), .B1(n712), .B2(n1351), .ZN(n1496) );
  OAI221_X1 U1534 ( .B1(n13), .B2(n715), .C1(n237), .C2(n718), .A(n1497), .ZN(
        n1492) );
  AOI22_X1 U1535 ( .A1(n721), .A2(n1179), .B1(n724), .B2(n1212), .ZN(n1497) );
  OAI221_X1 U1536 ( .B1(n14), .B2(n727), .C1(n238), .C2(n730), .A(n1498), .ZN(
        n1491) );
  AOI22_X1 U1537 ( .A1(n733), .A2(n1249), .B1(n736), .B2(n1282), .ZN(n1498) );
  NAND2_X1 U1538 ( .A1(n1499), .A2(n1500), .ZN(OUT2[7]) );
  NOR4_X1 U1539 ( .A1(n1501), .A2(n1502), .A3(n1503), .A4(n1504), .ZN(n1500)
         );
  OAI221_X1 U1540 ( .B1(n15), .B2(n643), .C1(n239), .C2(n646), .A(n1505), .ZN(
        n1504) );
  AOI22_X1 U1541 ( .A1(n649), .A2(n932), .B1(n652), .B2(n898), .ZN(n1505) );
  OAI221_X1 U1542 ( .B1(n16), .B2(n655), .C1(n240), .C2(n658), .A(n1506), .ZN(
        n1503) );
  AOI22_X1 U1543 ( .A1(n661), .A2(n1005), .B1(n664), .B2(n972), .ZN(n1506) );
  OAI221_X1 U1544 ( .B1(n17), .B2(n667), .C1(n241), .C2(n670), .A(n1507), .ZN(
        n1502) );
  AOI22_X1 U1545 ( .A1(n673), .A2(n1074), .B1(n676), .B2(n1041), .ZN(n1507) );
  OAI221_X1 U1546 ( .B1(n18), .B2(n679), .C1(n242), .C2(n682), .A(n1508), .ZN(
        n1501) );
  AOI22_X1 U1547 ( .A1(n685), .A2(n1143), .B1(n688), .B2(n1110), .ZN(n1508) );
  NOR4_X1 U1548 ( .A1(n1509), .A2(n1510), .A3(n1511), .A4(n1512), .ZN(n1499)
         );
  OAI221_X1 U1549 ( .B1(n3772), .B2(n691), .C1(n3773), .C2(n694), .A(n1513), 
        .ZN(n1512) );
  AOI22_X1 U1550 ( .A1(n697), .A2(n3774), .B1(n700), .B2(n3775), .ZN(n1513) );
  OAI221_X1 U1551 ( .B1(n19), .B2(n703), .C1(n243), .C2(n706), .A(n1514), .ZN(
        n1511) );
  AOI22_X1 U1552 ( .A1(n709), .A2(n1319), .B1(n712), .B2(n1352), .ZN(n1514) );
  OAI221_X1 U1553 ( .B1(n20), .B2(n715), .C1(n244), .C2(n718), .A(n1515), .ZN(
        n1510) );
  AOI22_X1 U1554 ( .A1(n721), .A2(n1180), .B1(n724), .B2(n1213), .ZN(n1515) );
  OAI221_X1 U1555 ( .B1(n21), .B2(n727), .C1(n245), .C2(n730), .A(n1516), .ZN(
        n1509) );
  AOI22_X1 U1556 ( .A1(n733), .A2(n1250), .B1(n736), .B2(n1283), .ZN(n1516) );
  NAND2_X1 U1557 ( .A1(n1517), .A2(n1518), .ZN(OUT2[6]) );
  NOR4_X1 U1558 ( .A1(n1519), .A2(n1520), .A3(n1521), .A4(n1522), .ZN(n1518)
         );
  OAI221_X1 U1559 ( .B1(n22), .B2(n643), .C1(n246), .C2(n646), .A(n1523), .ZN(
        n1522) );
  AOI22_X1 U1560 ( .A1(n649), .A2(n933), .B1(n652), .B2(n899), .ZN(n1523) );
  OAI221_X1 U1561 ( .B1(n23), .B2(n655), .C1(n247), .C2(n658), .A(n1524), .ZN(
        n1521) );
  AOI22_X1 U1562 ( .A1(n661), .A2(n1006), .B1(n664), .B2(n973), .ZN(n1524) );
  OAI221_X1 U1563 ( .B1(n24), .B2(n667), .C1(n248), .C2(n670), .A(n1525), .ZN(
        n1520) );
  AOI22_X1 U1564 ( .A1(n673), .A2(n1075), .B1(n676), .B2(n1042), .ZN(n1525) );
  OAI221_X1 U1565 ( .B1(n25), .B2(n679), .C1(n249), .C2(n682), .A(n1526), .ZN(
        n1519) );
  AOI22_X1 U1566 ( .A1(n685), .A2(n1144), .B1(n688), .B2(n1111), .ZN(n1526) );
  NOR4_X1 U1567 ( .A1(n1527), .A2(n1528), .A3(n1529), .A4(n1530), .ZN(n1517)
         );
  OAI221_X1 U1568 ( .B1(n3790), .B2(n691), .C1(n3791), .C2(n694), .A(n1531), 
        .ZN(n1530) );
  AOI22_X1 U1569 ( .A1(n697), .A2(n3792), .B1(n700), .B2(n3793), .ZN(n1531) );
  OAI221_X1 U1570 ( .B1(n26), .B2(n703), .C1(n250), .C2(n706), .A(n1532), .ZN(
        n1529) );
  AOI22_X1 U1571 ( .A1(n709), .A2(n1320), .B1(n712), .B2(n1353), .ZN(n1532) );
  OAI221_X1 U1572 ( .B1(n27), .B2(n715), .C1(n251), .C2(n718), .A(n1533), .ZN(
        n1528) );
  AOI22_X1 U1573 ( .A1(n721), .A2(n1181), .B1(n724), .B2(n1214), .ZN(n1533) );
  OAI221_X1 U1574 ( .B1(n28), .B2(n727), .C1(n252), .C2(n730), .A(n1534), .ZN(
        n1527) );
  AOI22_X1 U1575 ( .A1(n733), .A2(n1251), .B1(n736), .B2(n1284), .ZN(n1534) );
  NAND2_X1 U1576 ( .A1(n1535), .A2(n1536), .ZN(OUT2[5]) );
  NOR4_X1 U1577 ( .A1(n1537), .A2(n1538), .A3(n1539), .A4(n1540), .ZN(n1536)
         );
  OAI221_X1 U1578 ( .B1(n29), .B2(n643), .C1(n253), .C2(n646), .A(n1541), .ZN(
        n1540) );
  AOI22_X1 U1579 ( .A1(n649), .A2(n934), .B1(n652), .B2(n900), .ZN(n1541) );
  OAI221_X1 U1580 ( .B1(n30), .B2(n655), .C1(n254), .C2(n658), .A(n1542), .ZN(
        n1539) );
  AOI22_X1 U1581 ( .A1(n661), .A2(n1007), .B1(n664), .B2(n974), .ZN(n1542) );
  OAI221_X1 U1582 ( .B1(n31), .B2(n667), .C1(n255), .C2(n670), .A(n1543), .ZN(
        n1538) );
  AOI22_X1 U1583 ( .A1(n673), .A2(n1076), .B1(n676), .B2(n1043), .ZN(n1543) );
  OAI221_X1 U1584 ( .B1(n32), .B2(n679), .C1(n256), .C2(n682), .A(n1544), .ZN(
        n1537) );
  AOI22_X1 U1585 ( .A1(n685), .A2(n1145), .B1(n688), .B2(n1112), .ZN(n1544) );
  NOR4_X1 U1586 ( .A1(n1545), .A2(n1546), .A3(n1547), .A4(n1548), .ZN(n1535)
         );
  OAI221_X1 U1587 ( .B1(n3808), .B2(n691), .C1(n3809), .C2(n694), .A(n1549), 
        .ZN(n1548) );
  AOI22_X1 U1588 ( .A1(n697), .A2(n3810), .B1(n700), .B2(n3811), .ZN(n1549) );
  OAI221_X1 U1589 ( .B1(n33), .B2(n703), .C1(n257), .C2(n706), .A(n1550), .ZN(
        n1547) );
  AOI22_X1 U1590 ( .A1(n709), .A2(n1321), .B1(n712), .B2(n1354), .ZN(n1550) );
  OAI221_X1 U1591 ( .B1(n34), .B2(n715), .C1(n258), .C2(n718), .A(n1551), .ZN(
        n1546) );
  AOI22_X1 U1592 ( .A1(n721), .A2(n1182), .B1(n724), .B2(n1215), .ZN(n1551) );
  OAI221_X1 U1593 ( .B1(n35), .B2(n727), .C1(n259), .C2(n730), .A(n1552), .ZN(
        n1545) );
  AOI22_X1 U1594 ( .A1(n733), .A2(n1252), .B1(n736), .B2(n1285), .ZN(n1552) );
  NAND2_X1 U1595 ( .A1(n1553), .A2(n1554), .ZN(OUT2[4]) );
  NOR4_X1 U1596 ( .A1(n1555), .A2(n1556), .A3(n1557), .A4(n1558), .ZN(n1554)
         );
  OAI221_X1 U1597 ( .B1(n36), .B2(n643), .C1(n260), .C2(n646), .A(n1559), .ZN(
        n1558) );
  AOI22_X1 U1598 ( .A1(n649), .A2(n935), .B1(n652), .B2(n901), .ZN(n1559) );
  OAI221_X1 U1599 ( .B1(n37), .B2(n655), .C1(n261), .C2(n658), .A(n1560), .ZN(
        n1557) );
  AOI22_X1 U1600 ( .A1(n661), .A2(n1008), .B1(n664), .B2(n975), .ZN(n1560) );
  OAI221_X1 U1601 ( .B1(n38), .B2(n667), .C1(n262), .C2(n670), .A(n1561), .ZN(
        n1556) );
  AOI22_X1 U1602 ( .A1(n673), .A2(n1077), .B1(n676), .B2(n1044), .ZN(n1561) );
  OAI221_X1 U1603 ( .B1(n39), .B2(n679), .C1(n263), .C2(n682), .A(n1562), .ZN(
        n1555) );
  AOI22_X1 U1604 ( .A1(n685), .A2(n1146), .B1(n688), .B2(n1113), .ZN(n1562) );
  NOR4_X1 U1605 ( .A1(n1563), .A2(n1564), .A3(n1565), .A4(n1566), .ZN(n1553)
         );
  OAI221_X1 U1606 ( .B1(n3826), .B2(n691), .C1(n3827), .C2(n694), .A(n1567), 
        .ZN(n1566) );
  AOI22_X1 U1607 ( .A1(n697), .A2(n3828), .B1(n700), .B2(n3829), .ZN(n1567) );
  OAI221_X1 U1608 ( .B1(n40), .B2(n703), .C1(n264), .C2(n706), .A(n1568), .ZN(
        n1565) );
  AOI22_X1 U1609 ( .A1(n709), .A2(n1322), .B1(n712), .B2(n1355), .ZN(n1568) );
  OAI221_X1 U1610 ( .B1(n41), .B2(n715), .C1(n265), .C2(n718), .A(n1569), .ZN(
        n1564) );
  AOI22_X1 U1611 ( .A1(n721), .A2(n1183), .B1(n724), .B2(n1216), .ZN(n1569) );
  OAI221_X1 U1612 ( .B1(n42), .B2(n727), .C1(n266), .C2(n730), .A(n1570), .ZN(
        n1563) );
  AOI22_X1 U1613 ( .A1(n733), .A2(n1253), .B1(n736), .B2(n1286), .ZN(n1570) );
  NAND2_X1 U1614 ( .A1(n1571), .A2(n1572), .ZN(OUT2[3]) );
  NOR4_X1 U1615 ( .A1(n1573), .A2(n1574), .A3(n1575), .A4(n1576), .ZN(n1572)
         );
  OAI221_X1 U1616 ( .B1(n43), .B2(n643), .C1(n267), .C2(n646), .A(n1577), .ZN(
        n1576) );
  AOI22_X1 U1617 ( .A1(n649), .A2(n936), .B1(n652), .B2(n902), .ZN(n1577) );
  OAI221_X1 U1618 ( .B1(n44), .B2(n655), .C1(n268), .C2(n658), .A(n1578), .ZN(
        n1575) );
  AOI22_X1 U1619 ( .A1(n661), .A2(n1009), .B1(n664), .B2(n976), .ZN(n1578) );
  OAI221_X1 U1620 ( .B1(n45), .B2(n667), .C1(n269), .C2(n670), .A(n1579), .ZN(
        n1574) );
  AOI22_X1 U1621 ( .A1(n673), .A2(n1078), .B1(n676), .B2(n1045), .ZN(n1579) );
  OAI221_X1 U1622 ( .B1(n46), .B2(n679), .C1(n270), .C2(n682), .A(n1580), .ZN(
        n1573) );
  AOI22_X1 U1623 ( .A1(n685), .A2(n1147), .B1(n688), .B2(n1114), .ZN(n1580) );
  NOR4_X1 U1624 ( .A1(n1581), .A2(n1582), .A3(n1583), .A4(n1584), .ZN(n1571)
         );
  OAI221_X1 U1625 ( .B1(n3844), .B2(n691), .C1(n3845), .C2(n694), .A(n1585), 
        .ZN(n1584) );
  AOI22_X1 U1626 ( .A1(n697), .A2(n3846), .B1(n700), .B2(n3847), .ZN(n1585) );
  OAI221_X1 U1627 ( .B1(n47), .B2(n703), .C1(n271), .C2(n706), .A(n1586), .ZN(
        n1583) );
  AOI22_X1 U1628 ( .A1(n709), .A2(n1323), .B1(n712), .B2(n1356), .ZN(n1586) );
  OAI221_X1 U1629 ( .B1(n48), .B2(n715), .C1(n272), .C2(n718), .A(n1587), .ZN(
        n1582) );
  AOI22_X1 U1630 ( .A1(n721), .A2(n1184), .B1(n724), .B2(n1217), .ZN(n1587) );
  OAI221_X1 U1631 ( .B1(n49), .B2(n727), .C1(n273), .C2(n730), .A(n1588), .ZN(
        n1581) );
  AOI22_X1 U1632 ( .A1(n733), .A2(n1254), .B1(n736), .B2(n1287), .ZN(n1588) );
  NAND2_X1 U1633 ( .A1(n1589), .A2(n1590), .ZN(OUT2[31]) );
  NOR4_X1 U1634 ( .A1(n1591), .A2(n1592), .A3(n1593), .A4(n1594), .ZN(n1590)
         );
  OAI221_X1 U1635 ( .B1(n50), .B2(n643), .C1(n274), .C2(n646), .A(n1595), .ZN(
        n1594) );
  AOI22_X1 U1636 ( .A1(n649), .A2(n907), .B1(n652), .B2(n873), .ZN(n1595) );
  OAI221_X1 U1637 ( .B1(n51), .B2(n655), .C1(n275), .C2(n658), .A(n1596), .ZN(
        n1593) );
  AOI22_X1 U1638 ( .A1(n661), .A2(n980), .B1(n664), .B2(n947), .ZN(n1596) );
  OAI221_X1 U1639 ( .B1(n52), .B2(n667), .C1(n276), .C2(n670), .A(n1597), .ZN(
        n1592) );
  AOI22_X1 U1640 ( .A1(n673), .A2(n1049), .B1(n676), .B2(n1016), .ZN(n1597) );
  OAI221_X1 U1641 ( .B1(n53), .B2(n679), .C1(n277), .C2(n682), .A(n1598), .ZN(
        n1591) );
  AOI22_X1 U1642 ( .A1(n685), .A2(n1118), .B1(n688), .B2(n1085), .ZN(n1598) );
  NOR4_X1 U1643 ( .A1(n1599), .A2(n1600), .A3(n1601), .A4(n1602), .ZN(n1589)
         );
  OAI221_X1 U1644 ( .B1(n3862), .B2(n691), .C1(n3863), .C2(n694), .A(n1603), 
        .ZN(n1602) );
  AOI22_X1 U1645 ( .A1(n697), .A2(n3864), .B1(n700), .B2(n3865), .ZN(n1603) );
  OAI221_X1 U1646 ( .B1(n54), .B2(n703), .C1(n278), .C2(n706), .A(n1604), .ZN(
        n1601) );
  AOI22_X1 U1647 ( .A1(n709), .A2(n1294), .B1(n712), .B2(n1327), .ZN(n1604) );
  OAI221_X1 U1648 ( .B1(n55), .B2(n715), .C1(n279), .C2(n718), .A(n1605), .ZN(
        n1600) );
  AOI22_X1 U1649 ( .A1(n721), .A2(n1155), .B1(n724), .B2(n1188), .ZN(n1605) );
  OAI221_X1 U1650 ( .B1(n56), .B2(n727), .C1(n280), .C2(n730), .A(n1606), .ZN(
        n1599) );
  AOI22_X1 U1651 ( .A1(n733), .A2(n1225), .B1(n736), .B2(n1258), .ZN(n1606) );
  NAND2_X1 U1652 ( .A1(n1607), .A2(n1608), .ZN(OUT2[30]) );
  NOR4_X1 U1653 ( .A1(n1609), .A2(n1610), .A3(n1611), .A4(n1612), .ZN(n1608)
         );
  OAI221_X1 U1654 ( .B1(n57), .B2(n642), .C1(n281), .C2(n645), .A(n1613), .ZN(
        n1612) );
  AOI22_X1 U1655 ( .A1(n648), .A2(n909), .B1(n651), .B2(n875), .ZN(n1613) );
  OAI221_X1 U1656 ( .B1(n58), .B2(n654), .C1(n282), .C2(n657), .A(n1614), .ZN(
        n1611) );
  AOI22_X1 U1657 ( .A1(n660), .A2(n982), .B1(n663), .B2(n949), .ZN(n1614) );
  OAI221_X1 U1658 ( .B1(n59), .B2(n666), .C1(n283), .C2(n669), .A(n1615), .ZN(
        n1610) );
  AOI22_X1 U1659 ( .A1(n672), .A2(n1051), .B1(n675), .B2(n1018), .ZN(n1615) );
  OAI221_X1 U1660 ( .B1(n60), .B2(n678), .C1(n284), .C2(n681), .A(n1616), .ZN(
        n1609) );
  AOI22_X1 U1661 ( .A1(n684), .A2(n1120), .B1(n687), .B2(n1087), .ZN(n1616) );
  NOR4_X1 U1662 ( .A1(n1617), .A2(n1618), .A3(n1619), .A4(n1620), .ZN(n1607)
         );
  OAI221_X1 U1663 ( .B1(n3880), .B2(n690), .C1(n3881), .C2(n693), .A(n1621), 
        .ZN(n1620) );
  AOI22_X1 U1664 ( .A1(n696), .A2(n3882), .B1(n699), .B2(n3883), .ZN(n1621) );
  OAI221_X1 U1665 ( .B1(n61), .B2(n702), .C1(n285), .C2(n705), .A(n1622), .ZN(
        n1619) );
  AOI22_X1 U1666 ( .A1(n708), .A2(n1296), .B1(n711), .B2(n1329), .ZN(n1622) );
  OAI221_X1 U1667 ( .B1(n62), .B2(n714), .C1(n286), .C2(n717), .A(n1623), .ZN(
        n1618) );
  AOI22_X1 U1668 ( .A1(n720), .A2(n1157), .B1(n723), .B2(n1190), .ZN(n1623) );
  OAI221_X1 U1669 ( .B1(n63), .B2(n726), .C1(n287), .C2(n729), .A(n1624), .ZN(
        n1617) );
  AOI22_X1 U1670 ( .A1(n732), .A2(n1227), .B1(n735), .B2(n1260), .ZN(n1624) );
  NAND2_X1 U1671 ( .A1(n1625), .A2(n1626), .ZN(OUT2[2]) );
  NOR4_X1 U1672 ( .A1(n1627), .A2(n1628), .A3(n1629), .A4(n1630), .ZN(n1626)
         );
  OAI221_X1 U1673 ( .B1(n64), .B2(n642), .C1(n288), .C2(n645), .A(n1631), .ZN(
        n1630) );
  AOI22_X1 U1674 ( .A1(n648), .A2(n937), .B1(n651), .B2(n903), .ZN(n1631) );
  OAI221_X1 U1675 ( .B1(n65), .B2(n654), .C1(n289), .C2(n657), .A(n1632), .ZN(
        n1629) );
  AOI22_X1 U1676 ( .A1(n660), .A2(n1010), .B1(n663), .B2(n977), .ZN(n1632) );
  OAI221_X1 U1677 ( .B1(n66), .B2(n666), .C1(n290), .C2(n669), .A(n1633), .ZN(
        n1628) );
  AOI22_X1 U1678 ( .A1(n672), .A2(n1079), .B1(n675), .B2(n1046), .ZN(n1633) );
  OAI221_X1 U1679 ( .B1(n67), .B2(n678), .C1(n291), .C2(n681), .A(n1634), .ZN(
        n1627) );
  AOI22_X1 U1680 ( .A1(n684), .A2(n1148), .B1(n687), .B2(n1115), .ZN(n1634) );
  NOR4_X1 U1681 ( .A1(n1635), .A2(n1636), .A3(n1637), .A4(n1638), .ZN(n1625)
         );
  OAI221_X1 U1682 ( .B1(n3898), .B2(n690), .C1(n3899), .C2(n693), .A(n1639), 
        .ZN(n1638) );
  AOI22_X1 U1683 ( .A1(n696), .A2(n3900), .B1(n699), .B2(n3901), .ZN(n1639) );
  OAI221_X1 U1684 ( .B1(n68), .B2(n702), .C1(n292), .C2(n705), .A(n1640), .ZN(
        n1637) );
  AOI22_X1 U1685 ( .A1(n708), .A2(n1324), .B1(n711), .B2(n1357), .ZN(n1640) );
  OAI221_X1 U1686 ( .B1(n69), .B2(n714), .C1(n293), .C2(n717), .A(n1641), .ZN(
        n1636) );
  AOI22_X1 U1687 ( .A1(n720), .A2(n1185), .B1(n723), .B2(n1218), .ZN(n1641) );
  OAI221_X1 U1688 ( .B1(n70), .B2(n726), .C1(n294), .C2(n729), .A(n1642), .ZN(
        n1635) );
  AOI22_X1 U1689 ( .A1(n732), .A2(n1255), .B1(n735), .B2(n1288), .ZN(n1642) );
  NAND2_X1 U1690 ( .A1(n1643), .A2(n1644), .ZN(OUT2[29]) );
  NOR4_X1 U1691 ( .A1(n1645), .A2(n1646), .A3(n1647), .A4(n1648), .ZN(n1644)
         );
  OAI221_X1 U1692 ( .B1(n71), .B2(n642), .C1(n295), .C2(n645), .A(n1649), .ZN(
        n1648) );
  AOI22_X1 U1693 ( .A1(n648), .A2(n910), .B1(n651), .B2(n876), .ZN(n1649) );
  OAI221_X1 U1694 ( .B1(n72), .B2(n654), .C1(n296), .C2(n657), .A(n1650), .ZN(
        n1647) );
  AOI22_X1 U1695 ( .A1(n660), .A2(n983), .B1(n663), .B2(n950), .ZN(n1650) );
  OAI221_X1 U1696 ( .B1(n73), .B2(n666), .C1(n297), .C2(n669), .A(n1651), .ZN(
        n1646) );
  AOI22_X1 U1697 ( .A1(n672), .A2(n1052), .B1(n675), .B2(n1019), .ZN(n1651) );
  OAI221_X1 U1698 ( .B1(n74), .B2(n678), .C1(n298), .C2(n681), .A(n1652), .ZN(
        n1645) );
  AOI22_X1 U1699 ( .A1(n684), .A2(n1121), .B1(n687), .B2(n1088), .ZN(n1652) );
  NOR4_X1 U1700 ( .A1(n1653), .A2(n1654), .A3(n1655), .A4(n1656), .ZN(n1643)
         );
  OAI221_X1 U1701 ( .B1(n3916), .B2(n690), .C1(n3917), .C2(n693), .A(n1657), 
        .ZN(n1656) );
  AOI22_X1 U1702 ( .A1(n696), .A2(n3918), .B1(n699), .B2(n3919), .ZN(n1657) );
  OAI221_X1 U1703 ( .B1(n75), .B2(n702), .C1(n299), .C2(n705), .A(n1658), .ZN(
        n1655) );
  AOI22_X1 U1704 ( .A1(n708), .A2(n1297), .B1(n711), .B2(n1330), .ZN(n1658) );
  OAI221_X1 U1705 ( .B1(n76), .B2(n714), .C1(n300), .C2(n717), .A(n1659), .ZN(
        n1654) );
  AOI22_X1 U1706 ( .A1(n720), .A2(n1158), .B1(n723), .B2(n1191), .ZN(n1659) );
  OAI221_X1 U1707 ( .B1(n77), .B2(n726), .C1(n301), .C2(n729), .A(n1660), .ZN(
        n1653) );
  AOI22_X1 U1708 ( .A1(n732), .A2(n1228), .B1(n735), .B2(n1261), .ZN(n1660) );
  NAND2_X1 U1709 ( .A1(n1661), .A2(n1662), .ZN(OUT2[28]) );
  NOR4_X1 U1710 ( .A1(n1663), .A2(n1664), .A3(n1665), .A4(n1666), .ZN(n1662)
         );
  OAI221_X1 U1711 ( .B1(n78), .B2(n642), .C1(n302), .C2(n645), .A(n1667), .ZN(
        n1666) );
  AOI22_X1 U1712 ( .A1(n648), .A2(n911), .B1(n651), .B2(n877), .ZN(n1667) );
  OAI221_X1 U1713 ( .B1(n79), .B2(n654), .C1(n303), .C2(n657), .A(n1668), .ZN(
        n1665) );
  AOI22_X1 U1714 ( .A1(n660), .A2(n984), .B1(n663), .B2(n951), .ZN(n1668) );
  OAI221_X1 U1715 ( .B1(n80), .B2(n666), .C1(n304), .C2(n669), .A(n1669), .ZN(
        n1664) );
  AOI22_X1 U1716 ( .A1(n672), .A2(n1053), .B1(n675), .B2(n1020), .ZN(n1669) );
  OAI221_X1 U1717 ( .B1(n81), .B2(n678), .C1(n305), .C2(n681), .A(n1670), .ZN(
        n1663) );
  AOI22_X1 U1718 ( .A1(n684), .A2(n1122), .B1(n687), .B2(n1089), .ZN(n1670) );
  NOR4_X1 U1719 ( .A1(n1671), .A2(n1672), .A3(n1673), .A4(n1674), .ZN(n1661)
         );
  OAI221_X1 U1720 ( .B1(n3934), .B2(n690), .C1(n3935), .C2(n693), .A(n1675), 
        .ZN(n1674) );
  AOI22_X1 U1721 ( .A1(n696), .A2(n3936), .B1(n699), .B2(n3937), .ZN(n1675) );
  OAI221_X1 U1722 ( .B1(n82), .B2(n702), .C1(n306), .C2(n705), .A(n1676), .ZN(
        n1673) );
  AOI22_X1 U1723 ( .A1(n708), .A2(n1298), .B1(n711), .B2(n1331), .ZN(n1676) );
  OAI221_X1 U1724 ( .B1(n83), .B2(n714), .C1(n307), .C2(n717), .A(n1677), .ZN(
        n1672) );
  AOI22_X1 U1725 ( .A1(n720), .A2(n1159), .B1(n723), .B2(n1192), .ZN(n1677) );
  OAI221_X1 U1726 ( .B1(n84), .B2(n726), .C1(n308), .C2(n729), .A(n1678), .ZN(
        n1671) );
  AOI22_X1 U1727 ( .A1(n732), .A2(n1229), .B1(n735), .B2(n1262), .ZN(n1678) );
  NAND2_X1 U1728 ( .A1(n1679), .A2(n1680), .ZN(OUT2[27]) );
  NOR4_X1 U1729 ( .A1(n1681), .A2(n1682), .A3(n1683), .A4(n1684), .ZN(n1680)
         );
  OAI221_X1 U1730 ( .B1(n85), .B2(n642), .C1(n309), .C2(n645), .A(n1685), .ZN(
        n1684) );
  AOI22_X1 U1731 ( .A1(n648), .A2(n912), .B1(n651), .B2(n878), .ZN(n1685) );
  OAI221_X1 U1732 ( .B1(n86), .B2(n654), .C1(n310), .C2(n657), .A(n1686), .ZN(
        n1683) );
  AOI22_X1 U1733 ( .A1(n660), .A2(n985), .B1(n663), .B2(n952), .ZN(n1686) );
  OAI221_X1 U1734 ( .B1(n87), .B2(n666), .C1(n311), .C2(n669), .A(n1687), .ZN(
        n1682) );
  AOI22_X1 U1735 ( .A1(n672), .A2(n1054), .B1(n675), .B2(n1021), .ZN(n1687) );
  OAI221_X1 U1736 ( .B1(n88), .B2(n678), .C1(n312), .C2(n681), .A(n1688), .ZN(
        n1681) );
  AOI22_X1 U1737 ( .A1(n684), .A2(n1123), .B1(n687), .B2(n1090), .ZN(n1688) );
  NOR4_X1 U1738 ( .A1(n1689), .A2(n1690), .A3(n1691), .A4(n1692), .ZN(n1679)
         );
  OAI221_X1 U1739 ( .B1(n3952), .B2(n690), .C1(n3953), .C2(n693), .A(n1693), 
        .ZN(n1692) );
  AOI22_X1 U1740 ( .A1(n696), .A2(n3954), .B1(n699), .B2(n3955), .ZN(n1693) );
  OAI221_X1 U1741 ( .B1(n89), .B2(n702), .C1(n313), .C2(n705), .A(n1694), .ZN(
        n1691) );
  AOI22_X1 U1742 ( .A1(n708), .A2(n1299), .B1(n711), .B2(n1332), .ZN(n1694) );
  OAI221_X1 U1743 ( .B1(n90), .B2(n714), .C1(n314), .C2(n717), .A(n1695), .ZN(
        n1690) );
  AOI22_X1 U1744 ( .A1(n720), .A2(n1160), .B1(n723), .B2(n1193), .ZN(n1695) );
  OAI221_X1 U1745 ( .B1(n91), .B2(n726), .C1(n315), .C2(n729), .A(n1696), .ZN(
        n1689) );
  AOI22_X1 U1746 ( .A1(n732), .A2(n1230), .B1(n735), .B2(n1263), .ZN(n1696) );
  NAND2_X1 U1747 ( .A1(n1697), .A2(n1698), .ZN(OUT2[26]) );
  NOR4_X1 U1748 ( .A1(n1699), .A2(n1700), .A3(n1701), .A4(n1702), .ZN(n1698)
         );
  OAI221_X1 U1749 ( .B1(n92), .B2(n642), .C1(n316), .C2(n645), .A(n1703), .ZN(
        n1702) );
  AOI22_X1 U1750 ( .A1(n648), .A2(n913), .B1(n651), .B2(n879), .ZN(n1703) );
  OAI221_X1 U1751 ( .B1(n93), .B2(n654), .C1(n317), .C2(n657), .A(n1704), .ZN(
        n1701) );
  AOI22_X1 U1752 ( .A1(n660), .A2(n986), .B1(n663), .B2(n953), .ZN(n1704) );
  OAI221_X1 U1753 ( .B1(n94), .B2(n666), .C1(n318), .C2(n669), .A(n1705), .ZN(
        n1700) );
  AOI22_X1 U1754 ( .A1(n672), .A2(n1055), .B1(n675), .B2(n1022), .ZN(n1705) );
  OAI221_X1 U1755 ( .B1(n95), .B2(n678), .C1(n319), .C2(n681), .A(n1706), .ZN(
        n1699) );
  AOI22_X1 U1756 ( .A1(n684), .A2(n1124), .B1(n687), .B2(n1091), .ZN(n1706) );
  NOR4_X1 U1757 ( .A1(n1707), .A2(n1708), .A3(n1709), .A4(n1710), .ZN(n1697)
         );
  OAI221_X1 U1758 ( .B1(n3970), .B2(n690), .C1(n3971), .C2(n693), .A(n1711), 
        .ZN(n1710) );
  AOI22_X1 U1759 ( .A1(n696), .A2(n3972), .B1(n699), .B2(n3973), .ZN(n1711) );
  OAI221_X1 U1760 ( .B1(n96), .B2(n702), .C1(n320), .C2(n705), .A(n1712), .ZN(
        n1709) );
  AOI22_X1 U1761 ( .A1(n708), .A2(n1300), .B1(n711), .B2(n1333), .ZN(n1712) );
  OAI221_X1 U1762 ( .B1(n97), .B2(n714), .C1(n321), .C2(n717), .A(n1713), .ZN(
        n1708) );
  AOI22_X1 U1763 ( .A1(n720), .A2(n1161), .B1(n723), .B2(n1194), .ZN(n1713) );
  OAI221_X1 U1764 ( .B1(n98), .B2(n726), .C1(n322), .C2(n729), .A(n1714), .ZN(
        n1707) );
  AOI22_X1 U1765 ( .A1(n732), .A2(n1231), .B1(n735), .B2(n1264), .ZN(n1714) );
  NAND2_X1 U1766 ( .A1(n1715), .A2(n1716), .ZN(OUT2[25]) );
  NOR4_X1 U1767 ( .A1(n1717), .A2(n1718), .A3(n1719), .A4(n1720), .ZN(n1716)
         );
  OAI221_X1 U1768 ( .B1(n99), .B2(n642), .C1(n323), .C2(n645), .A(n1721), .ZN(
        n1720) );
  AOI22_X1 U1769 ( .A1(n648), .A2(n914), .B1(n651), .B2(n880), .ZN(n1721) );
  OAI221_X1 U1770 ( .B1(n100), .B2(n654), .C1(n324), .C2(n657), .A(n1722), 
        .ZN(n1719) );
  AOI22_X1 U1771 ( .A1(n660), .A2(n987), .B1(n663), .B2(n954), .ZN(n1722) );
  OAI221_X1 U1772 ( .B1(n101), .B2(n666), .C1(n325), .C2(n669), .A(n1723), 
        .ZN(n1718) );
  AOI22_X1 U1773 ( .A1(n672), .A2(n1056), .B1(n675), .B2(n1023), .ZN(n1723) );
  OAI221_X1 U1774 ( .B1(n102), .B2(n678), .C1(n326), .C2(n681), .A(n1724), 
        .ZN(n1717) );
  AOI22_X1 U1775 ( .A1(n684), .A2(n1125), .B1(n687), .B2(n1092), .ZN(n1724) );
  NOR4_X1 U1776 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(n1715)
         );
  OAI221_X1 U1777 ( .B1(n3988), .B2(n690), .C1(n3989), .C2(n693), .A(n1729), 
        .ZN(n1728) );
  AOI22_X1 U1778 ( .A1(n696), .A2(n3990), .B1(n699), .B2(n3991), .ZN(n1729) );
  OAI221_X1 U1779 ( .B1(n103), .B2(n702), .C1(n327), .C2(n705), .A(n1730), 
        .ZN(n1727) );
  AOI22_X1 U1780 ( .A1(n708), .A2(n1301), .B1(n711), .B2(n1334), .ZN(n1730) );
  OAI221_X1 U1781 ( .B1(n104), .B2(n714), .C1(n328), .C2(n717), .A(n1731), 
        .ZN(n1726) );
  AOI22_X1 U1782 ( .A1(n720), .A2(n1162), .B1(n723), .B2(n1195), .ZN(n1731) );
  OAI221_X1 U1783 ( .B1(n105), .B2(n726), .C1(n329), .C2(n729), .A(n1732), 
        .ZN(n1725) );
  AOI22_X1 U1784 ( .A1(n732), .A2(n1232), .B1(n735), .B2(n1265), .ZN(n1732) );
  NAND2_X1 U1785 ( .A1(n1733), .A2(n1734), .ZN(OUT2[24]) );
  NOR4_X1 U1786 ( .A1(n1735), .A2(n1736), .A3(n1737), .A4(n1738), .ZN(n1734)
         );
  OAI221_X1 U1787 ( .B1(n106), .B2(n642), .C1(n330), .C2(n645), .A(n1739), 
        .ZN(n1738) );
  AOI22_X1 U1788 ( .A1(n648), .A2(n915), .B1(n651), .B2(n881), .ZN(n1739) );
  OAI221_X1 U1789 ( .B1(n107), .B2(n654), .C1(n331), .C2(n657), .A(n1740), 
        .ZN(n1737) );
  AOI22_X1 U1790 ( .A1(n660), .A2(n988), .B1(n663), .B2(n955), .ZN(n1740) );
  OAI221_X1 U1791 ( .B1(n108), .B2(n666), .C1(n332), .C2(n669), .A(n1741), 
        .ZN(n1736) );
  AOI22_X1 U1792 ( .A1(n672), .A2(n1057), .B1(n675), .B2(n1024), .ZN(n1741) );
  OAI221_X1 U1793 ( .B1(n109), .B2(n678), .C1(n333), .C2(n681), .A(n1742), 
        .ZN(n1735) );
  AOI22_X1 U1794 ( .A1(n684), .A2(n1126), .B1(n687), .B2(n1093), .ZN(n1742) );
  NOR4_X1 U1795 ( .A1(n1743), .A2(n1744), .A3(n1745), .A4(n1746), .ZN(n1733)
         );
  OAI221_X1 U1796 ( .B1(n4006), .B2(n690), .C1(n4007), .C2(n693), .A(n1747), 
        .ZN(n1746) );
  AOI22_X1 U1797 ( .A1(n696), .A2(n4008), .B1(n699), .B2(n4009), .ZN(n1747) );
  OAI221_X1 U1798 ( .B1(n110), .B2(n702), .C1(n334), .C2(n705), .A(n1748), 
        .ZN(n1745) );
  AOI22_X1 U1799 ( .A1(n708), .A2(n1302), .B1(n711), .B2(n1335), .ZN(n1748) );
  OAI221_X1 U1800 ( .B1(n111), .B2(n714), .C1(n335), .C2(n717), .A(n1749), 
        .ZN(n1744) );
  AOI22_X1 U1801 ( .A1(n720), .A2(n1163), .B1(n723), .B2(n1196), .ZN(n1749) );
  OAI221_X1 U1802 ( .B1(n112), .B2(n726), .C1(n336), .C2(n729), .A(n1750), 
        .ZN(n1743) );
  AOI22_X1 U1803 ( .A1(n732), .A2(n1233), .B1(n735), .B2(n1266), .ZN(n1750) );
  NAND2_X1 U1804 ( .A1(n1751), .A2(n1752), .ZN(OUT2[23]) );
  NOR4_X1 U1805 ( .A1(n1753), .A2(n1754), .A3(n1755), .A4(n1756), .ZN(n1752)
         );
  OAI221_X1 U1806 ( .B1(n113), .B2(n642), .C1(n337), .C2(n645), .A(n1757), 
        .ZN(n1756) );
  AOI22_X1 U1807 ( .A1(n648), .A2(n916), .B1(n651), .B2(n882), .ZN(n1757) );
  OAI221_X1 U1808 ( .B1(n114), .B2(n654), .C1(n338), .C2(n657), .A(n1758), 
        .ZN(n1755) );
  AOI22_X1 U1809 ( .A1(n660), .A2(n989), .B1(n663), .B2(n956), .ZN(n1758) );
  OAI221_X1 U1810 ( .B1(n115), .B2(n666), .C1(n339), .C2(n669), .A(n1759), 
        .ZN(n1754) );
  AOI22_X1 U1811 ( .A1(n672), .A2(n1058), .B1(n675), .B2(n1025), .ZN(n1759) );
  OAI221_X1 U1812 ( .B1(n116), .B2(n678), .C1(n340), .C2(n681), .A(n1760), 
        .ZN(n1753) );
  AOI22_X1 U1813 ( .A1(n684), .A2(n1127), .B1(n687), .B2(n1094), .ZN(n1760) );
  NOR4_X1 U1814 ( .A1(n1761), .A2(n1762), .A3(n1763), .A4(n1764), .ZN(n1751)
         );
  OAI221_X1 U1815 ( .B1(n4024), .B2(n690), .C1(n4025), .C2(n693), .A(n1765), 
        .ZN(n1764) );
  AOI22_X1 U1816 ( .A1(n696), .A2(n4026), .B1(n699), .B2(n4027), .ZN(n1765) );
  OAI221_X1 U1817 ( .B1(n117), .B2(n702), .C1(n341), .C2(n705), .A(n1766), 
        .ZN(n1763) );
  AOI22_X1 U1818 ( .A1(n708), .A2(n1303), .B1(n711), .B2(n1336), .ZN(n1766) );
  OAI221_X1 U1819 ( .B1(n118), .B2(n714), .C1(n342), .C2(n717), .A(n1767), 
        .ZN(n1762) );
  AOI22_X1 U1820 ( .A1(n720), .A2(n1164), .B1(n723), .B2(n1197), .ZN(n1767) );
  OAI221_X1 U1821 ( .B1(n119), .B2(n726), .C1(n343), .C2(n729), .A(n1768), 
        .ZN(n1761) );
  AOI22_X1 U1822 ( .A1(n732), .A2(n1234), .B1(n735), .B2(n1267), .ZN(n1768) );
  NAND2_X1 U1823 ( .A1(n1769), .A2(n1770), .ZN(OUT2[22]) );
  NOR4_X1 U1824 ( .A1(n1771), .A2(n1772), .A3(n1773), .A4(n1774), .ZN(n1770)
         );
  OAI221_X1 U1825 ( .B1(n120), .B2(n642), .C1(n344), .C2(n645), .A(n1775), 
        .ZN(n1774) );
  AOI22_X1 U1826 ( .A1(n648), .A2(n917), .B1(n651), .B2(n883), .ZN(n1775) );
  OAI221_X1 U1827 ( .B1(n121), .B2(n654), .C1(n345), .C2(n657), .A(n1776), 
        .ZN(n1773) );
  AOI22_X1 U1828 ( .A1(n660), .A2(n990), .B1(n663), .B2(n957), .ZN(n1776) );
  OAI221_X1 U1829 ( .B1(n122), .B2(n666), .C1(n346), .C2(n669), .A(n1777), 
        .ZN(n1772) );
  AOI22_X1 U1830 ( .A1(n672), .A2(n1059), .B1(n675), .B2(n1026), .ZN(n1777) );
  OAI221_X1 U1831 ( .B1(n123), .B2(n678), .C1(n347), .C2(n681), .A(n1778), 
        .ZN(n1771) );
  AOI22_X1 U1832 ( .A1(n684), .A2(n1128), .B1(n687), .B2(n1095), .ZN(n1778) );
  NOR4_X1 U1833 ( .A1(n1779), .A2(n1780), .A3(n1781), .A4(n1782), .ZN(n1769)
         );
  OAI221_X1 U1834 ( .B1(n4042), .B2(n690), .C1(n4043), .C2(n693), .A(n1783), 
        .ZN(n1782) );
  AOI22_X1 U1835 ( .A1(n696), .A2(n4044), .B1(n699), .B2(n4045), .ZN(n1783) );
  OAI221_X1 U1836 ( .B1(n124), .B2(n702), .C1(n348), .C2(n705), .A(n1784), 
        .ZN(n1781) );
  AOI22_X1 U1837 ( .A1(n708), .A2(n1304), .B1(n711), .B2(n1337), .ZN(n1784) );
  OAI221_X1 U1838 ( .B1(n125), .B2(n714), .C1(n349), .C2(n717), .A(n1785), 
        .ZN(n1780) );
  AOI22_X1 U1839 ( .A1(n720), .A2(n1165), .B1(n723), .B2(n1198), .ZN(n1785) );
  OAI221_X1 U1840 ( .B1(n126), .B2(n726), .C1(n350), .C2(n729), .A(n1786), 
        .ZN(n1779) );
  AOI22_X1 U1841 ( .A1(n732), .A2(n1235), .B1(n735), .B2(n1268), .ZN(n1786) );
  NAND2_X1 U1842 ( .A1(n1787), .A2(n1788), .ZN(OUT2[21]) );
  NOR4_X1 U1843 ( .A1(n1789), .A2(n1790), .A3(n1791), .A4(n1792), .ZN(n1788)
         );
  OAI221_X1 U1844 ( .B1(n127), .B2(n642), .C1(n351), .C2(n645), .A(n1793), 
        .ZN(n1792) );
  AOI22_X1 U1845 ( .A1(n648), .A2(n918), .B1(n651), .B2(n884), .ZN(n1793) );
  OAI221_X1 U1846 ( .B1(n128), .B2(n654), .C1(n352), .C2(n657), .A(n1794), 
        .ZN(n1791) );
  AOI22_X1 U1847 ( .A1(n660), .A2(n991), .B1(n663), .B2(n958), .ZN(n1794) );
  OAI221_X1 U1848 ( .B1(n129), .B2(n666), .C1(n353), .C2(n669), .A(n1795), 
        .ZN(n1790) );
  AOI22_X1 U1849 ( .A1(n672), .A2(n1060), .B1(n675), .B2(n1027), .ZN(n1795) );
  OAI221_X1 U1850 ( .B1(n130), .B2(n678), .C1(n354), .C2(n681), .A(n1796), 
        .ZN(n1789) );
  AOI22_X1 U1851 ( .A1(n684), .A2(n1129), .B1(n687), .B2(n1096), .ZN(n1796) );
  NOR4_X1 U1852 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .ZN(n1787)
         );
  OAI221_X1 U1853 ( .B1(n4060), .B2(n690), .C1(n4061), .C2(n693), .A(n1801), 
        .ZN(n1800) );
  AOI22_X1 U1854 ( .A1(n696), .A2(n4062), .B1(n699), .B2(n4063), .ZN(n1801) );
  OAI221_X1 U1855 ( .B1(n131), .B2(n702), .C1(n355), .C2(n705), .A(n1802), 
        .ZN(n1799) );
  AOI22_X1 U1856 ( .A1(n708), .A2(n1305), .B1(n711), .B2(n1338), .ZN(n1802) );
  OAI221_X1 U1857 ( .B1(n132), .B2(n714), .C1(n356), .C2(n717), .A(n1803), 
        .ZN(n1798) );
  AOI22_X1 U1858 ( .A1(n720), .A2(n1166), .B1(n723), .B2(n1199), .ZN(n1803) );
  OAI221_X1 U1859 ( .B1(n133), .B2(n726), .C1(n357), .C2(n729), .A(n1804), 
        .ZN(n1797) );
  AOI22_X1 U1860 ( .A1(n732), .A2(n1236), .B1(n735), .B2(n1269), .ZN(n1804) );
  NAND2_X1 U1861 ( .A1(n1805), .A2(n1806), .ZN(OUT2[20]) );
  NOR4_X1 U1862 ( .A1(n1807), .A2(n1808), .A3(n1809), .A4(n1810), .ZN(n1806)
         );
  OAI221_X1 U1863 ( .B1(n134), .B2(n642), .C1(n358), .C2(n645), .A(n1811), 
        .ZN(n1810) );
  AOI22_X1 U1864 ( .A1(n648), .A2(n919), .B1(n651), .B2(n885), .ZN(n1811) );
  OAI221_X1 U1865 ( .B1(n135), .B2(n654), .C1(n359), .C2(n657), .A(n1812), 
        .ZN(n1809) );
  AOI22_X1 U1866 ( .A1(n660), .A2(n992), .B1(n663), .B2(n959), .ZN(n1812) );
  OAI221_X1 U1867 ( .B1(n136), .B2(n666), .C1(n360), .C2(n669), .A(n1813), 
        .ZN(n1808) );
  AOI22_X1 U1868 ( .A1(n672), .A2(n1061), .B1(n675), .B2(n1028), .ZN(n1813) );
  OAI221_X1 U1869 ( .B1(n137), .B2(n678), .C1(n361), .C2(n681), .A(n1814), 
        .ZN(n1807) );
  AOI22_X1 U1870 ( .A1(n684), .A2(n1130), .B1(n687), .B2(n1097), .ZN(n1814) );
  NOR4_X1 U1871 ( .A1(n1815), .A2(n1816), .A3(n1817), .A4(n1818), .ZN(n1805)
         );
  OAI221_X1 U1872 ( .B1(n4078), .B2(n690), .C1(n4079), .C2(n693), .A(n1819), 
        .ZN(n1818) );
  AOI22_X1 U1873 ( .A1(n696), .A2(n4080), .B1(n699), .B2(n4081), .ZN(n1819) );
  OAI221_X1 U1874 ( .B1(n138), .B2(n702), .C1(n362), .C2(n705), .A(n1820), 
        .ZN(n1817) );
  AOI22_X1 U1875 ( .A1(n708), .A2(n1306), .B1(n711), .B2(n1339), .ZN(n1820) );
  OAI221_X1 U1876 ( .B1(n139), .B2(n714), .C1(n363), .C2(n717), .A(n1821), 
        .ZN(n1816) );
  AOI22_X1 U1877 ( .A1(n720), .A2(n1167), .B1(n723), .B2(n1200), .ZN(n1821) );
  OAI221_X1 U1878 ( .B1(n140), .B2(n726), .C1(n364), .C2(n729), .A(n1822), 
        .ZN(n1815) );
  AOI22_X1 U1879 ( .A1(n732), .A2(n1237), .B1(n735), .B2(n1270), .ZN(n1822) );
  NAND2_X1 U1880 ( .A1(n1823), .A2(n1824), .ZN(OUT2[1]) );
  NOR4_X1 U1881 ( .A1(n1825), .A2(n1826), .A3(n1827), .A4(n1828), .ZN(n1824)
         );
  OAI221_X1 U1882 ( .B1(n141), .B2(n641), .C1(n365), .C2(n644), .A(n1829), 
        .ZN(n1828) );
  AOI22_X1 U1883 ( .A1(n647), .A2(n938), .B1(n650), .B2(n904), .ZN(n1829) );
  OAI221_X1 U1884 ( .B1(n142), .B2(n653), .C1(n366), .C2(n656), .A(n1830), 
        .ZN(n1827) );
  AOI22_X1 U1885 ( .A1(n659), .A2(n1011), .B1(n662), .B2(n978), .ZN(n1830) );
  OAI221_X1 U1886 ( .B1(n143), .B2(n665), .C1(n367), .C2(n668), .A(n1831), 
        .ZN(n1826) );
  AOI22_X1 U1887 ( .A1(n671), .A2(n1080), .B1(n674), .B2(n1047), .ZN(n1831) );
  OAI221_X1 U1888 ( .B1(n144), .B2(n677), .C1(n368), .C2(n680), .A(n1832), 
        .ZN(n1825) );
  AOI22_X1 U1889 ( .A1(n683), .A2(n1149), .B1(n686), .B2(n1116), .ZN(n1832) );
  NOR4_X1 U1890 ( .A1(n1833), .A2(n1834), .A3(n1835), .A4(n1836), .ZN(n1823)
         );
  OAI221_X1 U1891 ( .B1(n4096), .B2(n689), .C1(n4097), .C2(n692), .A(n1837), 
        .ZN(n1836) );
  AOI22_X1 U1892 ( .A1(n695), .A2(n4098), .B1(n698), .B2(n4099), .ZN(n1837) );
  OAI221_X1 U1893 ( .B1(n145), .B2(n701), .C1(n369), .C2(n704), .A(n1838), 
        .ZN(n1835) );
  AOI22_X1 U1894 ( .A1(n707), .A2(n1325), .B1(n710), .B2(n1358), .ZN(n1838) );
  OAI221_X1 U1895 ( .B1(n146), .B2(n713), .C1(n370), .C2(n716), .A(n1839), 
        .ZN(n1834) );
  AOI22_X1 U1896 ( .A1(n719), .A2(n1186), .B1(n722), .B2(n1219), .ZN(n1839) );
  OAI221_X1 U1897 ( .B1(n147), .B2(n725), .C1(n371), .C2(n728), .A(n1840), 
        .ZN(n1833) );
  AOI22_X1 U1898 ( .A1(n731), .A2(n1256), .B1(n734), .B2(n1289), .ZN(n1840) );
  NAND2_X1 U1899 ( .A1(n1841), .A2(n1842), .ZN(OUT2[19]) );
  NOR4_X1 U1900 ( .A1(n1843), .A2(n1844), .A3(n1845), .A4(n1846), .ZN(n1842)
         );
  OAI221_X1 U1901 ( .B1(n148), .B2(n641), .C1(n372), .C2(n644), .A(n1847), 
        .ZN(n1846) );
  AOI22_X1 U1902 ( .A1(n647), .A2(n920), .B1(n650), .B2(n886), .ZN(n1847) );
  OAI221_X1 U1903 ( .B1(n149), .B2(n653), .C1(n373), .C2(n656), .A(n1848), 
        .ZN(n1845) );
  AOI22_X1 U1904 ( .A1(n659), .A2(n993), .B1(n662), .B2(n960), .ZN(n1848) );
  OAI221_X1 U1905 ( .B1(n150), .B2(n665), .C1(n374), .C2(n668), .A(n1849), 
        .ZN(n1844) );
  AOI22_X1 U1906 ( .A1(n671), .A2(n1062), .B1(n674), .B2(n1029), .ZN(n1849) );
  OAI221_X1 U1907 ( .B1(n151), .B2(n677), .C1(n375), .C2(n680), .A(n1850), 
        .ZN(n1843) );
  AOI22_X1 U1908 ( .A1(n683), .A2(n1131), .B1(n686), .B2(n1098), .ZN(n1850) );
  NOR4_X1 U1909 ( .A1(n1851), .A2(n1852), .A3(n1853), .A4(n1854), .ZN(n1841)
         );
  OAI221_X1 U1910 ( .B1(n4114), .B2(n689), .C1(n4115), .C2(n692), .A(n1855), 
        .ZN(n1854) );
  AOI22_X1 U1911 ( .A1(n695), .A2(n4116), .B1(n698), .B2(n4117), .ZN(n1855) );
  OAI221_X1 U1912 ( .B1(n152), .B2(n701), .C1(n376), .C2(n704), .A(n1856), 
        .ZN(n1853) );
  AOI22_X1 U1913 ( .A1(n707), .A2(n1307), .B1(n710), .B2(n1340), .ZN(n1856) );
  OAI221_X1 U1914 ( .B1(n153), .B2(n713), .C1(n377), .C2(n716), .A(n1857), 
        .ZN(n1852) );
  AOI22_X1 U1915 ( .A1(n719), .A2(n1168), .B1(n722), .B2(n1201), .ZN(n1857) );
  OAI221_X1 U1916 ( .B1(n154), .B2(n725), .C1(n378), .C2(n728), .A(n1858), 
        .ZN(n1851) );
  AOI22_X1 U1917 ( .A1(n731), .A2(n1238), .B1(n734), .B2(n1271), .ZN(n1858) );
  NAND2_X1 U1918 ( .A1(n1859), .A2(n1860), .ZN(OUT2[18]) );
  NOR4_X1 U1919 ( .A1(n1861), .A2(n1862), .A3(n1863), .A4(n1864), .ZN(n1860)
         );
  OAI221_X1 U1920 ( .B1(n155), .B2(n641), .C1(n379), .C2(n644), .A(n1865), 
        .ZN(n1864) );
  AOI22_X1 U1921 ( .A1(n647), .A2(n921), .B1(n650), .B2(n887), .ZN(n1865) );
  OAI221_X1 U1922 ( .B1(n156), .B2(n653), .C1(n380), .C2(n656), .A(n1866), 
        .ZN(n1863) );
  AOI22_X1 U1923 ( .A1(n659), .A2(n994), .B1(n662), .B2(n961), .ZN(n1866) );
  OAI221_X1 U1924 ( .B1(n157), .B2(n665), .C1(n381), .C2(n668), .A(n1867), 
        .ZN(n1862) );
  AOI22_X1 U1925 ( .A1(n671), .A2(n1063), .B1(n674), .B2(n1030), .ZN(n1867) );
  OAI221_X1 U1926 ( .B1(n158), .B2(n677), .C1(n382), .C2(n680), .A(n1868), 
        .ZN(n1861) );
  AOI22_X1 U1927 ( .A1(n683), .A2(n1132), .B1(n686), .B2(n1099), .ZN(n1868) );
  NOR4_X1 U1928 ( .A1(n1869), .A2(n1870), .A3(n1871), .A4(n1872), .ZN(n1859)
         );
  OAI221_X1 U1929 ( .B1(n4132), .B2(n689), .C1(n4133), .C2(n692), .A(n1873), 
        .ZN(n1872) );
  AOI22_X1 U1930 ( .A1(n695), .A2(n4134), .B1(n698), .B2(n4135), .ZN(n1873) );
  OAI221_X1 U1931 ( .B1(n159), .B2(n701), .C1(n383), .C2(n704), .A(n1874), 
        .ZN(n1871) );
  AOI22_X1 U1932 ( .A1(n707), .A2(n1308), .B1(n710), .B2(n1341), .ZN(n1874) );
  OAI221_X1 U1933 ( .B1(n160), .B2(n713), .C1(n384), .C2(n716), .A(n1875), 
        .ZN(n1870) );
  AOI22_X1 U1934 ( .A1(n719), .A2(n1169), .B1(n722), .B2(n1202), .ZN(n1875) );
  OAI221_X1 U1935 ( .B1(n161), .B2(n725), .C1(n385), .C2(n728), .A(n1876), 
        .ZN(n1869) );
  AOI22_X1 U1936 ( .A1(n731), .A2(n1239), .B1(n734), .B2(n1272), .ZN(n1876) );
  NAND2_X1 U1937 ( .A1(n1877), .A2(n1878), .ZN(OUT2[17]) );
  NOR4_X1 U1938 ( .A1(n1879), .A2(n1880), .A3(n1881), .A4(n1882), .ZN(n1878)
         );
  OAI221_X1 U1939 ( .B1(n162), .B2(n641), .C1(n386), .C2(n644), .A(n1883), 
        .ZN(n1882) );
  AOI22_X1 U1940 ( .A1(n647), .A2(n922), .B1(n650), .B2(n888), .ZN(n1883) );
  OAI221_X1 U1941 ( .B1(n163), .B2(n653), .C1(n387), .C2(n656), .A(n1884), 
        .ZN(n1881) );
  AOI22_X1 U1942 ( .A1(n659), .A2(n995), .B1(n662), .B2(n962), .ZN(n1884) );
  OAI221_X1 U1943 ( .B1(n164), .B2(n665), .C1(n388), .C2(n668), .A(n1885), 
        .ZN(n1880) );
  AOI22_X1 U1944 ( .A1(n671), .A2(n1064), .B1(n674), .B2(n1031), .ZN(n1885) );
  OAI221_X1 U1945 ( .B1(n165), .B2(n677), .C1(n389), .C2(n680), .A(n1886), 
        .ZN(n1879) );
  AOI22_X1 U1946 ( .A1(n683), .A2(n1133), .B1(n686), .B2(n1100), .ZN(n1886) );
  NOR4_X1 U1947 ( .A1(n1887), .A2(n1888), .A3(n1889), .A4(n1890), .ZN(n1877)
         );
  OAI221_X1 U1948 ( .B1(n4150), .B2(n689), .C1(n4151), .C2(n692), .A(n1891), 
        .ZN(n1890) );
  AOI22_X1 U1949 ( .A1(n695), .A2(n4152), .B1(n698), .B2(n4153), .ZN(n1891) );
  OAI221_X1 U1950 ( .B1(n166), .B2(n701), .C1(n390), .C2(n704), .A(n1892), 
        .ZN(n1889) );
  AOI22_X1 U1951 ( .A1(n707), .A2(n1309), .B1(n710), .B2(n1342), .ZN(n1892) );
  OAI221_X1 U1952 ( .B1(n167), .B2(n713), .C1(n391), .C2(n716), .A(n1893), 
        .ZN(n1888) );
  AOI22_X1 U1953 ( .A1(n719), .A2(n1170), .B1(n722), .B2(n1203), .ZN(n1893) );
  OAI221_X1 U1954 ( .B1(n168), .B2(n725), .C1(n392), .C2(n728), .A(n1894), 
        .ZN(n1887) );
  AOI22_X1 U1955 ( .A1(n731), .A2(n1240), .B1(n734), .B2(n1273), .ZN(n1894) );
  NAND2_X1 U1956 ( .A1(n1895), .A2(n1896), .ZN(OUT2[16]) );
  NOR4_X1 U1957 ( .A1(n1897), .A2(n1898), .A3(n1899), .A4(n1900), .ZN(n1896)
         );
  OAI221_X1 U1958 ( .B1(n169), .B2(n641), .C1(n393), .C2(n644), .A(n1901), 
        .ZN(n1900) );
  AOI22_X1 U1959 ( .A1(n647), .A2(n923), .B1(n650), .B2(n889), .ZN(n1901) );
  OAI221_X1 U1960 ( .B1(n170), .B2(n653), .C1(n394), .C2(n656), .A(n1902), 
        .ZN(n1899) );
  AOI22_X1 U1961 ( .A1(n659), .A2(n996), .B1(n662), .B2(n963), .ZN(n1902) );
  OAI221_X1 U1962 ( .B1(n171), .B2(n665), .C1(n395), .C2(n668), .A(n1903), 
        .ZN(n1898) );
  AOI22_X1 U1963 ( .A1(n671), .A2(n1065), .B1(n674), .B2(n1032), .ZN(n1903) );
  OAI221_X1 U1964 ( .B1(n172), .B2(n677), .C1(n396), .C2(n680), .A(n1904), 
        .ZN(n1897) );
  AOI22_X1 U1965 ( .A1(n683), .A2(n1134), .B1(n686), .B2(n1101), .ZN(n1904) );
  NOR4_X1 U1966 ( .A1(n1905), .A2(n1906), .A3(n1907), .A4(n1908), .ZN(n1895)
         );
  OAI221_X1 U1967 ( .B1(n4168), .B2(n689), .C1(n4169), .C2(n692), .A(n1909), 
        .ZN(n1908) );
  AOI22_X1 U1968 ( .A1(n695), .A2(n4170), .B1(n698), .B2(n4171), .ZN(n1909) );
  OAI221_X1 U1969 ( .B1(n173), .B2(n701), .C1(n397), .C2(n704), .A(n1910), 
        .ZN(n1907) );
  AOI22_X1 U1970 ( .A1(n707), .A2(n1310), .B1(n710), .B2(n1343), .ZN(n1910) );
  OAI221_X1 U1971 ( .B1(n174), .B2(n713), .C1(n398), .C2(n716), .A(n1911), 
        .ZN(n1906) );
  AOI22_X1 U1972 ( .A1(n719), .A2(n1171), .B1(n722), .B2(n1204), .ZN(n1911) );
  OAI221_X1 U1973 ( .B1(n175), .B2(n725), .C1(n399), .C2(n728), .A(n1912), 
        .ZN(n1905) );
  AOI22_X1 U1974 ( .A1(n731), .A2(n1241), .B1(n734), .B2(n1274), .ZN(n1912) );
  NAND2_X1 U1975 ( .A1(n1913), .A2(n1914), .ZN(OUT2[15]) );
  NOR4_X1 U1976 ( .A1(n1915), .A2(n1916), .A3(n1917), .A4(n1918), .ZN(n1914)
         );
  OAI221_X1 U1977 ( .B1(n176), .B2(n641), .C1(n400), .C2(n644), .A(n1919), 
        .ZN(n1918) );
  AOI22_X1 U1978 ( .A1(n647), .A2(n924), .B1(n650), .B2(n890), .ZN(n1919) );
  OAI221_X1 U1979 ( .B1(n177), .B2(n653), .C1(n401), .C2(n656), .A(n1920), 
        .ZN(n1917) );
  AOI22_X1 U1980 ( .A1(n659), .A2(n997), .B1(n662), .B2(n964), .ZN(n1920) );
  OAI221_X1 U1981 ( .B1(n178), .B2(n665), .C1(n402), .C2(n668), .A(n1921), 
        .ZN(n1916) );
  AOI22_X1 U1982 ( .A1(n671), .A2(n1066), .B1(n674), .B2(n1033), .ZN(n1921) );
  OAI221_X1 U1983 ( .B1(n179), .B2(n677), .C1(n403), .C2(n680), .A(n1922), 
        .ZN(n1915) );
  AOI22_X1 U1984 ( .A1(n683), .A2(n1135), .B1(n686), .B2(n1102), .ZN(n1922) );
  NOR4_X1 U1985 ( .A1(n1923), .A2(n1924), .A3(n1925), .A4(n1926), .ZN(n1913)
         );
  OAI221_X1 U1986 ( .B1(n4186), .B2(n689), .C1(n4187), .C2(n692), .A(n1927), 
        .ZN(n1926) );
  AOI22_X1 U1987 ( .A1(n695), .A2(n4188), .B1(n698), .B2(n4189), .ZN(n1927) );
  OAI221_X1 U1988 ( .B1(n180), .B2(n701), .C1(n404), .C2(n704), .A(n1928), 
        .ZN(n1925) );
  AOI22_X1 U1989 ( .A1(n707), .A2(n1311), .B1(n710), .B2(n1344), .ZN(n1928) );
  OAI221_X1 U1990 ( .B1(n181), .B2(n713), .C1(n405), .C2(n716), .A(n1929), 
        .ZN(n1924) );
  AOI22_X1 U1991 ( .A1(n719), .A2(n1172), .B1(n722), .B2(n1205), .ZN(n1929) );
  OAI221_X1 U1992 ( .B1(n182), .B2(n725), .C1(n406), .C2(n728), .A(n1930), 
        .ZN(n1923) );
  AOI22_X1 U1993 ( .A1(n731), .A2(n1242), .B1(n734), .B2(n1275), .ZN(n1930) );
  NAND2_X1 U1994 ( .A1(n1931), .A2(n1932), .ZN(OUT2[14]) );
  NOR4_X1 U1995 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(n1932)
         );
  OAI221_X1 U1996 ( .B1(n183), .B2(n641), .C1(n407), .C2(n644), .A(n1937), 
        .ZN(n1936) );
  AOI22_X1 U1997 ( .A1(n647), .A2(n925), .B1(n650), .B2(n891), .ZN(n1937) );
  OAI221_X1 U1998 ( .B1(n184), .B2(n653), .C1(n408), .C2(n656), .A(n1938), 
        .ZN(n1935) );
  AOI22_X1 U1999 ( .A1(n659), .A2(n998), .B1(n662), .B2(n965), .ZN(n1938) );
  OAI221_X1 U2000 ( .B1(n185), .B2(n665), .C1(n409), .C2(n668), .A(n1939), 
        .ZN(n1934) );
  AOI22_X1 U2001 ( .A1(n671), .A2(n1067), .B1(n674), .B2(n1034), .ZN(n1939) );
  OAI221_X1 U2002 ( .B1(n186), .B2(n677), .C1(n410), .C2(n680), .A(n1940), 
        .ZN(n1933) );
  AOI22_X1 U2003 ( .A1(n683), .A2(n1136), .B1(n686), .B2(n1103), .ZN(n1940) );
  NOR4_X1 U2004 ( .A1(n1941), .A2(n1942), .A3(n1943), .A4(n1944), .ZN(n1931)
         );
  OAI221_X1 U2005 ( .B1(n4204), .B2(n689), .C1(n4205), .C2(n692), .A(n1945), 
        .ZN(n1944) );
  AOI22_X1 U2006 ( .A1(n695), .A2(n4206), .B1(n698), .B2(n4207), .ZN(n1945) );
  OAI221_X1 U2007 ( .B1(n187), .B2(n701), .C1(n411), .C2(n704), .A(n1946), 
        .ZN(n1943) );
  AOI22_X1 U2008 ( .A1(n707), .A2(n1312), .B1(n710), .B2(n1345), .ZN(n1946) );
  OAI221_X1 U2009 ( .B1(n188), .B2(n713), .C1(n412), .C2(n716), .A(n1947), 
        .ZN(n1942) );
  AOI22_X1 U2010 ( .A1(n719), .A2(n1173), .B1(n722), .B2(n1206), .ZN(n1947) );
  OAI221_X1 U2011 ( .B1(n189), .B2(n725), .C1(n413), .C2(n728), .A(n1948), 
        .ZN(n1941) );
  AOI22_X1 U2012 ( .A1(n731), .A2(n1243), .B1(n734), .B2(n1276), .ZN(n1948) );
  NAND2_X1 U2013 ( .A1(n1949), .A2(n1950), .ZN(OUT2[13]) );
  NOR4_X1 U2014 ( .A1(n1951), .A2(n1952), .A3(n1953), .A4(n1954), .ZN(n1950)
         );
  OAI221_X1 U2015 ( .B1(n190), .B2(n641), .C1(n414), .C2(n644), .A(n1955), 
        .ZN(n1954) );
  AOI22_X1 U2016 ( .A1(n647), .A2(n926), .B1(n650), .B2(n892), .ZN(n1955) );
  OAI221_X1 U2017 ( .B1(n191), .B2(n653), .C1(n415), .C2(n656), .A(n1956), 
        .ZN(n1953) );
  AOI22_X1 U2018 ( .A1(n659), .A2(n999), .B1(n662), .B2(n966), .ZN(n1956) );
  OAI221_X1 U2019 ( .B1(n192), .B2(n665), .C1(n416), .C2(n668), .A(n1957), 
        .ZN(n1952) );
  AOI22_X1 U2020 ( .A1(n671), .A2(n1068), .B1(n674), .B2(n1035), .ZN(n1957) );
  OAI221_X1 U2021 ( .B1(n193), .B2(n677), .C1(n417), .C2(n680), .A(n1958), 
        .ZN(n1951) );
  AOI22_X1 U2022 ( .A1(n683), .A2(n1137), .B1(n686), .B2(n1104), .ZN(n1958) );
  NOR4_X1 U2023 ( .A1(n1959), .A2(n1960), .A3(n1961), .A4(n1962), .ZN(n1949)
         );
  OAI221_X1 U2024 ( .B1(n4222), .B2(n689), .C1(n4223), .C2(n692), .A(n1963), 
        .ZN(n1962) );
  AOI22_X1 U2025 ( .A1(n695), .A2(n4224), .B1(n698), .B2(n4225), .ZN(n1963) );
  OAI221_X1 U2026 ( .B1(n194), .B2(n701), .C1(n418), .C2(n704), .A(n1964), 
        .ZN(n1961) );
  AOI22_X1 U2027 ( .A1(n707), .A2(n1313), .B1(n710), .B2(n1346), .ZN(n1964) );
  OAI221_X1 U2028 ( .B1(n195), .B2(n713), .C1(n419), .C2(n716), .A(n1965), 
        .ZN(n1960) );
  AOI22_X1 U2029 ( .A1(n719), .A2(n1174), .B1(n722), .B2(n1207), .ZN(n1965) );
  OAI221_X1 U2030 ( .B1(n196), .B2(n725), .C1(n420), .C2(n728), .A(n1966), 
        .ZN(n1959) );
  AOI22_X1 U2031 ( .A1(n731), .A2(n1244), .B1(n734), .B2(n1277), .ZN(n1966) );
  NAND2_X1 U2032 ( .A1(n1967), .A2(n1968), .ZN(OUT2[12]) );
  NOR4_X1 U2033 ( .A1(n1969), .A2(n1970), .A3(n1971), .A4(n1972), .ZN(n1968)
         );
  OAI221_X1 U2034 ( .B1(n197), .B2(n641), .C1(n421), .C2(n644), .A(n1973), 
        .ZN(n1972) );
  AOI22_X1 U2035 ( .A1(n647), .A2(n927), .B1(n650), .B2(n893), .ZN(n1973) );
  OAI221_X1 U2036 ( .B1(n198), .B2(n653), .C1(n422), .C2(n656), .A(n1974), 
        .ZN(n1971) );
  AOI22_X1 U2037 ( .A1(n659), .A2(n1000), .B1(n662), .B2(n967), .ZN(n1974) );
  OAI221_X1 U2038 ( .B1(n199), .B2(n665), .C1(n423), .C2(n668), .A(n1975), 
        .ZN(n1970) );
  AOI22_X1 U2039 ( .A1(n671), .A2(n1069), .B1(n674), .B2(n1036), .ZN(n1975) );
  OAI221_X1 U2040 ( .B1(n200), .B2(n677), .C1(n424), .C2(n680), .A(n1976), 
        .ZN(n1969) );
  AOI22_X1 U2041 ( .A1(n683), .A2(n1138), .B1(n686), .B2(n1105), .ZN(n1976) );
  NOR4_X1 U2042 ( .A1(n1977), .A2(n1978), .A3(n1979), .A4(n1980), .ZN(n1967)
         );
  OAI221_X1 U2043 ( .B1(n4240), .B2(n689), .C1(n4241), .C2(n692), .A(n1981), 
        .ZN(n1980) );
  AOI22_X1 U2044 ( .A1(n695), .A2(n4242), .B1(n698), .B2(n4243), .ZN(n1981) );
  OAI221_X1 U2045 ( .B1(n201), .B2(n701), .C1(n425), .C2(n704), .A(n1982), 
        .ZN(n1979) );
  AOI22_X1 U2046 ( .A1(n707), .A2(n1314), .B1(n710), .B2(n1347), .ZN(n1982) );
  OAI221_X1 U2047 ( .B1(n202), .B2(n713), .C1(n426), .C2(n716), .A(n1983), 
        .ZN(n1978) );
  AOI22_X1 U2048 ( .A1(n719), .A2(n1175), .B1(n722), .B2(n1208), .ZN(n1983) );
  OAI221_X1 U2049 ( .B1(n203), .B2(n725), .C1(n427), .C2(n728), .A(n1984), 
        .ZN(n1977) );
  AOI22_X1 U2050 ( .A1(n731), .A2(n1245), .B1(n734), .B2(n1278), .ZN(n1984) );
  NAND2_X1 U2051 ( .A1(n1985), .A2(n1986), .ZN(OUT2[11]) );
  NOR4_X1 U2052 ( .A1(n1987), .A2(n1988), .A3(n1989), .A4(n1990), .ZN(n1986)
         );
  OAI221_X1 U2053 ( .B1(n204), .B2(n641), .C1(n428), .C2(n644), .A(n1991), 
        .ZN(n1990) );
  AOI22_X1 U2054 ( .A1(n647), .A2(n928), .B1(n650), .B2(n894), .ZN(n1991) );
  OAI221_X1 U2055 ( .B1(n205), .B2(n653), .C1(n429), .C2(n656), .A(n1992), 
        .ZN(n1989) );
  AOI22_X1 U2056 ( .A1(n659), .A2(n1001), .B1(n662), .B2(n968), .ZN(n1992) );
  OAI221_X1 U2057 ( .B1(n206), .B2(n665), .C1(n430), .C2(n668), .A(n1993), 
        .ZN(n1988) );
  AOI22_X1 U2058 ( .A1(n671), .A2(n1070), .B1(n674), .B2(n1037), .ZN(n1993) );
  OAI221_X1 U2059 ( .B1(n207), .B2(n677), .C1(n431), .C2(n680), .A(n1994), 
        .ZN(n1987) );
  AOI22_X1 U2060 ( .A1(n683), .A2(n1139), .B1(n686), .B2(n1106), .ZN(n1994) );
  NOR4_X1 U2061 ( .A1(n1995), .A2(n1996), .A3(n1997), .A4(n1998), .ZN(n1985)
         );
  OAI221_X1 U2062 ( .B1(n4258), .B2(n689), .C1(n4259), .C2(n692), .A(n1999), 
        .ZN(n1998) );
  AOI22_X1 U2063 ( .A1(n695), .A2(n4260), .B1(n698), .B2(n4261), .ZN(n1999) );
  OAI221_X1 U2064 ( .B1(n208), .B2(n701), .C1(n432), .C2(n704), .A(n2000), 
        .ZN(n1997) );
  AOI22_X1 U2065 ( .A1(n707), .A2(n1315), .B1(n710), .B2(n1348), .ZN(n2000) );
  OAI221_X1 U2066 ( .B1(n209), .B2(n713), .C1(n433), .C2(n716), .A(n2001), 
        .ZN(n1996) );
  AOI22_X1 U2067 ( .A1(n719), .A2(n1176), .B1(n722), .B2(n1209), .ZN(n2001) );
  OAI221_X1 U2068 ( .B1(n210), .B2(n725), .C1(n434), .C2(n728), .A(n2002), 
        .ZN(n1995) );
  AOI22_X1 U2069 ( .A1(n731), .A2(n1246), .B1(n734), .B2(n1279), .ZN(n2002) );
  NAND2_X1 U2070 ( .A1(n2003), .A2(n2004), .ZN(OUT2[10]) );
  NOR4_X1 U2071 ( .A1(n2005), .A2(n2006), .A3(n2007), .A4(n2008), .ZN(n2004)
         );
  OAI221_X1 U2072 ( .B1(n211), .B2(n641), .C1(n435), .C2(n644), .A(n2009), 
        .ZN(n2008) );
  AOI22_X1 U2073 ( .A1(n647), .A2(n929), .B1(n650), .B2(n895), .ZN(n2009) );
  OAI221_X1 U2074 ( .B1(n212), .B2(n653), .C1(n436), .C2(n656), .A(n2010), 
        .ZN(n2007) );
  AOI22_X1 U2075 ( .A1(n659), .A2(n1002), .B1(n662), .B2(n969), .ZN(n2010) );
  OAI221_X1 U2076 ( .B1(n213), .B2(n665), .C1(n437), .C2(n668), .A(n2011), 
        .ZN(n2006) );
  AOI22_X1 U2077 ( .A1(n671), .A2(n1071), .B1(n674), .B2(n1038), .ZN(n2011) );
  OAI221_X1 U2078 ( .B1(n214), .B2(n677), .C1(n438), .C2(n680), .A(n2012), 
        .ZN(n2005) );
  AOI22_X1 U2079 ( .A1(n683), .A2(n1140), .B1(n686), .B2(n1107), .ZN(n2012) );
  NOR4_X1 U2080 ( .A1(n2013), .A2(n2014), .A3(n2015), .A4(n2016), .ZN(n2003)
         );
  OAI221_X1 U2081 ( .B1(n4276), .B2(n689), .C1(n4277), .C2(n692), .A(n2017), 
        .ZN(n2016) );
  AOI22_X1 U2082 ( .A1(n695), .A2(n4278), .B1(n698), .B2(n4279), .ZN(n2017) );
  OAI221_X1 U2083 ( .B1(n215), .B2(n701), .C1(n439), .C2(n704), .A(n2018), 
        .ZN(n2015) );
  AOI22_X1 U2084 ( .A1(n707), .A2(n1316), .B1(n710), .B2(n1349), .ZN(n2018) );
  OAI221_X1 U2085 ( .B1(n216), .B2(n713), .C1(n440), .C2(n716), .A(n2019), 
        .ZN(n2014) );
  AOI22_X1 U2086 ( .A1(n719), .A2(n1177), .B1(n722), .B2(n1210), .ZN(n2019) );
  OAI221_X1 U2087 ( .B1(n217), .B2(n725), .C1(n441), .C2(n728), .A(n2020), 
        .ZN(n2013) );
  AOI22_X1 U2088 ( .A1(n731), .A2(n1247), .B1(n734), .B2(n1280), .ZN(n2020) );
  NAND2_X1 U2089 ( .A1(n2021), .A2(n2022), .ZN(OUT2[0]) );
  NOR4_X1 U2090 ( .A1(n2023), .A2(n2024), .A3(n2025), .A4(n2026), .ZN(n2022)
         );
  OAI221_X1 U2091 ( .B1(n218), .B2(n641), .C1(n442), .C2(n644), .A(n2027), 
        .ZN(n2026) );
  AOI22_X1 U2092 ( .A1(n647), .A2(n939), .B1(n650), .B2(n905), .ZN(n2027) );
  AND2_X1 U2093 ( .A1(n2028), .A2(n2029), .ZN(n1441) );
  AND2_X1 U2094 ( .A1(n2030), .A2(n2029), .ZN(n1440) );
  NAND2_X1 U2095 ( .A1(n2028), .A2(n2031), .ZN(n1438) );
  NAND2_X1 U2096 ( .A1(n2030), .A2(n2031), .ZN(n1437) );
  OAI221_X1 U2097 ( .B1(n219), .B2(n653), .C1(n443), .C2(n656), .A(n2032), 
        .ZN(n2025) );
  AOI22_X1 U2098 ( .A1(n659), .A2(n1012), .B1(n662), .B2(n979), .ZN(n2032) );
  AND2_X1 U2099 ( .A1(n2028), .A2(n2033), .ZN(n1446) );
  AND2_X1 U2100 ( .A1(n2030), .A2(n2033), .ZN(n1445) );
  NAND2_X1 U2101 ( .A1(n2028), .A2(n2034), .ZN(n1443) );
  NOR3_X1 U2102 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n2028) );
  NAND2_X1 U2103 ( .A1(n2030), .A2(n2034), .ZN(n1442) );
  NOR3_X1 U2104 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n2035), .ZN(n2030) );
  OAI221_X1 U2105 ( .B1(n220), .B2(n665), .C1(n444), .C2(n668), .A(n2036), 
        .ZN(n2024) );
  AOI22_X1 U2106 ( .A1(n671), .A2(n1081), .B1(n674), .B2(n1048), .ZN(n2036) );
  AND2_X1 U2107 ( .A1(n2029), .A2(n2037), .ZN(n1451) );
  AND2_X1 U2108 ( .A1(n2029), .A2(n2038), .ZN(n1450) );
  NAND2_X1 U2109 ( .A1(n2031), .A2(n2037), .ZN(n1448) );
  NAND2_X1 U2110 ( .A1(n2031), .A2(n2038), .ZN(n1447) );
  OAI221_X1 U2111 ( .B1(n221), .B2(n677), .C1(n445), .C2(n680), .A(n2039), 
        .ZN(n2023) );
  AOI22_X1 U2112 ( .A1(n683), .A2(n1150), .B1(n686), .B2(n1117), .ZN(n2039) );
  AND2_X1 U2113 ( .A1(n2037), .A2(n2033), .ZN(n1456) );
  AND2_X1 U2114 ( .A1(n2038), .A2(n2033), .ZN(n1455) );
  NAND2_X1 U2115 ( .A1(n2034), .A2(n2037), .ZN(n1453) );
  NOR3_X1 U2116 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n2040), .ZN(n2037) );
  NAND2_X1 U2117 ( .A1(n2034), .A2(n2038), .ZN(n1452) );
  NOR3_X1 U2118 ( .A1(n2035), .A2(ADD_RD2[4]), .A3(n2040), .ZN(n2038) );
  NOR4_X1 U2119 ( .A1(n2041), .A2(n2042), .A3(n2043), .A4(n2044), .ZN(n2021)
         );
  OAI221_X1 U2120 ( .B1(n4294), .B2(n689), .C1(n4295), .C2(n692), .A(n2045), 
        .ZN(n2044) );
  AOI22_X1 U2121 ( .A1(n695), .A2(n4296), .B1(n698), .B2(n4297), .ZN(n2045) );
  AND2_X1 U2122 ( .A1(n2046), .A2(n2033), .ZN(n1465) );
  AND2_X1 U2123 ( .A1(n2047), .A2(n2033), .ZN(n1464) );
  NAND2_X1 U2124 ( .A1(n2047), .A2(n2034), .ZN(n1462) );
  NAND2_X1 U2125 ( .A1(n2046), .A2(n2034), .ZN(n1461) );
  OAI221_X1 U2126 ( .B1(n222), .B2(n701), .C1(n446), .C2(n704), .A(n2048), 
        .ZN(n2043) );
  AOI22_X1 U2127 ( .A1(n707), .A2(n1326), .B1(n710), .B2(n1359), .ZN(n2048) );
  AND2_X1 U2128 ( .A1(n2047), .A2(n2029), .ZN(n1470) );
  AND2_X1 U2129 ( .A1(n2046), .A2(n2029), .ZN(n1469) );
  NAND2_X1 U2130 ( .A1(n2046), .A2(n2031), .ZN(n1467) );
  NOR3_X1 U2131 ( .A1(n2040), .A2(ADD_RD2[0]), .A3(n2049), .ZN(n2046) );
  NAND2_X1 U2132 ( .A1(n2047), .A2(n2031), .ZN(n1466) );
  NOR3_X1 U2133 ( .A1(n2040), .A2(n2035), .A3(n2049), .ZN(n2047) );
  INV_X1 U2134 ( .A(ADD_RD2[3]), .ZN(n2040) );
  OAI221_X1 U2135 ( .B1(n223), .B2(n713), .C1(n447), .C2(n716), .A(n2050), 
        .ZN(n2042) );
  AOI22_X1 U2136 ( .A1(n719), .A2(n1187), .B1(n722), .B2(n1220), .ZN(n2050) );
  AND2_X1 U2137 ( .A1(n2051), .A2(n2029), .ZN(n1475) );
  AND2_X1 U2138 ( .A1(n2052), .A2(n2029), .ZN(n1474) );
  NOR3_X1 U2139 ( .A1(n2053), .A2(ADD_RD2[2]), .A3(n2054), .ZN(n2029) );
  NAND2_X1 U2140 ( .A1(n2051), .A2(n2031), .ZN(n1472) );
  NAND2_X1 U2141 ( .A1(n2052), .A2(n2031), .ZN(n1471) );
  OAI221_X1 U2142 ( .B1(n224), .B2(n725), .C1(n448), .C2(n728), .A(n2055), 
        .ZN(n2041) );
  AOI22_X1 U2143 ( .A1(n731), .A2(n1257), .B1(n734), .B2(n1290), .ZN(n2055) );
  AND2_X1 U2144 ( .A1(n2051), .A2(n2033), .ZN(n1480) );
  AND2_X1 U2145 ( .A1(n2052), .A2(n2033), .ZN(n1479) );
  NOR3_X1 U2146 ( .A1(n2056), .A2(n2053), .A3(n2054), .ZN(n2033) );
  NAND2_X1 U2147 ( .A1(n2051), .A2(n2034), .ZN(n1477) );
  NOR3_X1 U2148 ( .A1(n2035), .A2(ADD_RD2[3]), .A3(n2049), .ZN(n2051) );
  INV_X1 U2149 ( .A(ADD_RD2[0]), .ZN(n2035) );
  NAND2_X1 U2150 ( .A1(n2052), .A2(n2034), .ZN(n1476) );
  NOR3_X1 U2151 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n2049), .ZN(n2052) );
  NAND2_X1 U2152 ( .A1(n2057), .A2(n2058), .ZN(OUT1[9]) );
  NOR4_X1 U2153 ( .A1(n2059), .A2(n2060), .A3(n2061), .A4(n2062), .ZN(n2058)
         );
  OAI221_X1 U2154 ( .B1(n1), .B2(n739), .C1(n225), .C2(n742), .A(n2065), .ZN(
        n2062) );
  AOI22_X1 U2155 ( .A1(n745), .A2(n930), .B1(n748), .B2(n896), .ZN(n2065) );
  OAI221_X1 U2156 ( .B1(n2), .B2(n751), .C1(n226), .C2(n754), .A(n2070), .ZN(
        n2061) );
  AOI22_X1 U2157 ( .A1(n757), .A2(n1003), .B1(n760), .B2(n970), .ZN(n2070) );
  OAI221_X1 U2158 ( .B1(n3), .B2(n763), .C1(n227), .C2(n766), .A(n2075), .ZN(
        n2060) );
  AOI22_X1 U2159 ( .A1(n769), .A2(n1072), .B1(n772), .B2(n1039), .ZN(n2075) );
  OAI221_X1 U2160 ( .B1(n4), .B2(n775), .C1(n228), .C2(n778), .A(n2080), .ZN(
        n2059) );
  AOI22_X1 U2161 ( .A1(n781), .A2(n1141), .B1(n784), .B2(n1108), .ZN(n2080) );
  NOR4_X1 U2162 ( .A1(n2083), .A2(n2084), .A3(n2085), .A4(n2086), .ZN(n2057)
         );
  OAI221_X1 U2163 ( .B1(n3736), .B2(n787), .C1(n3737), .C2(n790), .A(n2089), 
        .ZN(n2086) );
  AOI22_X1 U2164 ( .A1(n793), .A2(n3738), .B1(n796), .B2(n3739), .ZN(n2089) );
  OAI221_X1 U2165 ( .B1(n5), .B2(n799), .C1(n229), .C2(n802), .A(n2094), .ZN(
        n2085) );
  AOI22_X1 U2166 ( .A1(n805), .A2(n1317), .B1(n808), .B2(n1350), .ZN(n2094) );
  OAI221_X1 U2167 ( .B1(n6), .B2(n811), .C1(n230), .C2(n814), .A(n2099), .ZN(
        n2084) );
  AOI22_X1 U2168 ( .A1(n817), .A2(n1178), .B1(n820), .B2(n1211), .ZN(n2099) );
  OAI221_X1 U2169 ( .B1(n7), .B2(n823), .C1(n231), .C2(n826), .A(n2104), .ZN(
        n2083) );
  AOI22_X1 U2170 ( .A1(n829), .A2(n1248), .B1(n832), .B2(n1281), .ZN(n2104) );
  NAND2_X1 U2171 ( .A1(n2107), .A2(n2108), .ZN(OUT1[8]) );
  NOR4_X1 U2172 ( .A1(n2109), .A2(n2110), .A3(n2111), .A4(n2112), .ZN(n2108)
         );
  OAI221_X1 U2173 ( .B1(n8), .B2(n739), .C1(n232), .C2(n742), .A(n2113), .ZN(
        n2112) );
  AOI22_X1 U2174 ( .A1(n745), .A2(n931), .B1(n748), .B2(n897), .ZN(n2113) );
  OAI221_X1 U2175 ( .B1(n9), .B2(n751), .C1(n233), .C2(n754), .A(n2114), .ZN(
        n2111) );
  AOI22_X1 U2176 ( .A1(n757), .A2(n1004), .B1(n760), .B2(n971), .ZN(n2114) );
  OAI221_X1 U2177 ( .B1(n10), .B2(n763), .C1(n234), .C2(n766), .A(n2115), .ZN(
        n2110) );
  AOI22_X1 U2178 ( .A1(n769), .A2(n1073), .B1(n772), .B2(n1040), .ZN(n2115) );
  OAI221_X1 U2179 ( .B1(n11), .B2(n775), .C1(n235), .C2(n778), .A(n2116), .ZN(
        n2109) );
  AOI22_X1 U2180 ( .A1(n781), .A2(n1142), .B1(n784), .B2(n1109), .ZN(n2116) );
  NOR4_X1 U2181 ( .A1(n2117), .A2(n2118), .A3(n2119), .A4(n2120), .ZN(n2107)
         );
  OAI221_X1 U2182 ( .B1(n3754), .B2(n787), .C1(n3755), .C2(n790), .A(n2121), 
        .ZN(n2120) );
  AOI22_X1 U2183 ( .A1(n793), .A2(n3756), .B1(n796), .B2(n3757), .ZN(n2121) );
  OAI221_X1 U2184 ( .B1(n12), .B2(n799), .C1(n236), .C2(n802), .A(n2122), .ZN(
        n2119) );
  AOI22_X1 U2185 ( .A1(n805), .A2(n1318), .B1(n808), .B2(n1351), .ZN(n2122) );
  OAI221_X1 U2186 ( .B1(n13), .B2(n811), .C1(n237), .C2(n814), .A(n2123), .ZN(
        n2118) );
  AOI22_X1 U2187 ( .A1(n817), .A2(n1179), .B1(n820), .B2(n1212), .ZN(n2123) );
  OAI221_X1 U2188 ( .B1(n14), .B2(n823), .C1(n238), .C2(n826), .A(n2124), .ZN(
        n2117) );
  AOI22_X1 U2189 ( .A1(n829), .A2(n1249), .B1(n832), .B2(n1282), .ZN(n2124) );
  NAND2_X1 U2190 ( .A1(n2125), .A2(n2126), .ZN(OUT1[7]) );
  NOR4_X1 U2191 ( .A1(n2127), .A2(n2128), .A3(n2129), .A4(n2130), .ZN(n2126)
         );
  OAI221_X1 U2192 ( .B1(n15), .B2(n739), .C1(n239), .C2(n742), .A(n2131), .ZN(
        n2130) );
  AOI22_X1 U2193 ( .A1(n745), .A2(n932), .B1(n748), .B2(n898), .ZN(n2131) );
  OAI221_X1 U2194 ( .B1(n16), .B2(n751), .C1(n240), .C2(n754), .A(n2132), .ZN(
        n2129) );
  AOI22_X1 U2195 ( .A1(n757), .A2(n1005), .B1(n760), .B2(n972), .ZN(n2132) );
  OAI221_X1 U2196 ( .B1(n17), .B2(n763), .C1(n241), .C2(n766), .A(n2133), .ZN(
        n2128) );
  AOI22_X1 U2197 ( .A1(n769), .A2(n1074), .B1(n772), .B2(n1041), .ZN(n2133) );
  OAI221_X1 U2198 ( .B1(n18), .B2(n775), .C1(n242), .C2(n778), .A(n2134), .ZN(
        n2127) );
  AOI22_X1 U2199 ( .A1(n781), .A2(n1143), .B1(n784), .B2(n1110), .ZN(n2134) );
  NOR4_X1 U2200 ( .A1(n2135), .A2(n2136), .A3(n2137), .A4(n2138), .ZN(n2125)
         );
  OAI221_X1 U2201 ( .B1(n3772), .B2(n787), .C1(n3773), .C2(n790), .A(n2139), 
        .ZN(n2138) );
  AOI22_X1 U2202 ( .A1(n793), .A2(n3774), .B1(n796), .B2(n3775), .ZN(n2139) );
  OAI221_X1 U2203 ( .B1(n19), .B2(n799), .C1(n243), .C2(n802), .A(n2140), .ZN(
        n2137) );
  AOI22_X1 U2204 ( .A1(n805), .A2(n1319), .B1(n808), .B2(n1352), .ZN(n2140) );
  OAI221_X1 U2205 ( .B1(n20), .B2(n811), .C1(n244), .C2(n814), .A(n2141), .ZN(
        n2136) );
  AOI22_X1 U2206 ( .A1(n817), .A2(n1180), .B1(n820), .B2(n1213), .ZN(n2141) );
  OAI221_X1 U2207 ( .B1(n21), .B2(n823), .C1(n245), .C2(n826), .A(n2142), .ZN(
        n2135) );
  AOI22_X1 U2208 ( .A1(n829), .A2(n1250), .B1(n832), .B2(n1283), .ZN(n2142) );
  NAND2_X1 U2209 ( .A1(n2143), .A2(n2144), .ZN(OUT1[6]) );
  NOR4_X1 U2210 ( .A1(n2145), .A2(n2146), .A3(n2147), .A4(n2148), .ZN(n2144)
         );
  OAI221_X1 U2211 ( .B1(n22), .B2(n739), .C1(n246), .C2(n742), .A(n2149), .ZN(
        n2148) );
  AOI22_X1 U2212 ( .A1(n745), .A2(n933), .B1(n748), .B2(n899), .ZN(n2149) );
  OAI221_X1 U2213 ( .B1(n23), .B2(n751), .C1(n247), .C2(n754), .A(n2150), .ZN(
        n2147) );
  AOI22_X1 U2214 ( .A1(n757), .A2(n1006), .B1(n760), .B2(n973), .ZN(n2150) );
  OAI221_X1 U2215 ( .B1(n24), .B2(n763), .C1(n248), .C2(n766), .A(n2151), .ZN(
        n2146) );
  AOI22_X1 U2216 ( .A1(n769), .A2(n1075), .B1(n772), .B2(n1042), .ZN(n2151) );
  OAI221_X1 U2217 ( .B1(n25), .B2(n775), .C1(n249), .C2(n778), .A(n2152), .ZN(
        n2145) );
  AOI22_X1 U2218 ( .A1(n781), .A2(n1144), .B1(n784), .B2(n1111), .ZN(n2152) );
  NOR4_X1 U2219 ( .A1(n2153), .A2(n2154), .A3(n2155), .A4(n2156), .ZN(n2143)
         );
  OAI221_X1 U2220 ( .B1(n3790), .B2(n787), .C1(n3791), .C2(n790), .A(n2157), 
        .ZN(n2156) );
  AOI22_X1 U2221 ( .A1(n793), .A2(n3792), .B1(n796), .B2(n3793), .ZN(n2157) );
  OAI221_X1 U2222 ( .B1(n26), .B2(n799), .C1(n250), .C2(n802), .A(n2158), .ZN(
        n2155) );
  AOI22_X1 U2223 ( .A1(n805), .A2(n1320), .B1(n808), .B2(n1353), .ZN(n2158) );
  OAI221_X1 U2224 ( .B1(n27), .B2(n811), .C1(n251), .C2(n814), .A(n2159), .ZN(
        n2154) );
  AOI22_X1 U2225 ( .A1(n817), .A2(n1181), .B1(n820), .B2(n1214), .ZN(n2159) );
  OAI221_X1 U2226 ( .B1(n28), .B2(n823), .C1(n252), .C2(n826), .A(n2160), .ZN(
        n2153) );
  AOI22_X1 U2227 ( .A1(n829), .A2(n1251), .B1(n832), .B2(n1284), .ZN(n2160) );
  NAND2_X1 U2228 ( .A1(n2161), .A2(n2162), .ZN(OUT1[5]) );
  NOR4_X1 U2229 ( .A1(n2163), .A2(n2164), .A3(n2165), .A4(n2166), .ZN(n2162)
         );
  OAI221_X1 U2230 ( .B1(n29), .B2(n739), .C1(n253), .C2(n742), .A(n2167), .ZN(
        n2166) );
  AOI22_X1 U2231 ( .A1(n745), .A2(n934), .B1(n748), .B2(n900), .ZN(n2167) );
  OAI221_X1 U2232 ( .B1(n30), .B2(n751), .C1(n254), .C2(n754), .A(n2168), .ZN(
        n2165) );
  AOI22_X1 U2233 ( .A1(n757), .A2(n1007), .B1(n760), .B2(n974), .ZN(n2168) );
  OAI221_X1 U2234 ( .B1(n31), .B2(n763), .C1(n255), .C2(n766), .A(n2169), .ZN(
        n2164) );
  AOI22_X1 U2235 ( .A1(n769), .A2(n1076), .B1(n772), .B2(n1043), .ZN(n2169) );
  OAI221_X1 U2236 ( .B1(n32), .B2(n775), .C1(n256), .C2(n778), .A(n2170), .ZN(
        n2163) );
  AOI22_X1 U2237 ( .A1(n781), .A2(n1145), .B1(n784), .B2(n1112), .ZN(n2170) );
  NOR4_X1 U2238 ( .A1(n2171), .A2(n2172), .A3(n2173), .A4(n2174), .ZN(n2161)
         );
  OAI221_X1 U2239 ( .B1(n3808), .B2(n787), .C1(n3809), .C2(n790), .A(n2175), 
        .ZN(n2174) );
  AOI22_X1 U2240 ( .A1(n793), .A2(n3810), .B1(n796), .B2(n3811), .ZN(n2175) );
  OAI221_X1 U2241 ( .B1(n33), .B2(n799), .C1(n257), .C2(n802), .A(n2176), .ZN(
        n2173) );
  AOI22_X1 U2242 ( .A1(n805), .A2(n1321), .B1(n808), .B2(n1354), .ZN(n2176) );
  OAI221_X1 U2243 ( .B1(n34), .B2(n811), .C1(n258), .C2(n814), .A(n2177), .ZN(
        n2172) );
  AOI22_X1 U2244 ( .A1(n817), .A2(n1182), .B1(n820), .B2(n1215), .ZN(n2177) );
  OAI221_X1 U2245 ( .B1(n35), .B2(n823), .C1(n259), .C2(n826), .A(n2178), .ZN(
        n2171) );
  AOI22_X1 U2246 ( .A1(n829), .A2(n1252), .B1(n832), .B2(n1285), .ZN(n2178) );
  NAND2_X1 U2247 ( .A1(n2179), .A2(n2180), .ZN(OUT1[4]) );
  NOR4_X1 U2248 ( .A1(n2181), .A2(n2182), .A3(n2183), .A4(n2184), .ZN(n2180)
         );
  OAI221_X1 U2249 ( .B1(n36), .B2(n739), .C1(n260), .C2(n742), .A(n2185), .ZN(
        n2184) );
  AOI22_X1 U2250 ( .A1(n745), .A2(n935), .B1(n748), .B2(n901), .ZN(n2185) );
  OAI221_X1 U2251 ( .B1(n37), .B2(n751), .C1(n261), .C2(n754), .A(n2186), .ZN(
        n2183) );
  AOI22_X1 U2252 ( .A1(n757), .A2(n1008), .B1(n760), .B2(n975), .ZN(n2186) );
  OAI221_X1 U2253 ( .B1(n38), .B2(n763), .C1(n262), .C2(n766), .A(n2187), .ZN(
        n2182) );
  AOI22_X1 U2254 ( .A1(n769), .A2(n1077), .B1(n772), .B2(n1044), .ZN(n2187) );
  OAI221_X1 U2255 ( .B1(n39), .B2(n775), .C1(n263), .C2(n778), .A(n2188), .ZN(
        n2181) );
  AOI22_X1 U2256 ( .A1(n781), .A2(n1146), .B1(n784), .B2(n1113), .ZN(n2188) );
  NOR4_X1 U2257 ( .A1(n2189), .A2(n2190), .A3(n2191), .A4(n2192), .ZN(n2179)
         );
  OAI221_X1 U2258 ( .B1(n3826), .B2(n787), .C1(n3827), .C2(n790), .A(n2193), 
        .ZN(n2192) );
  AOI22_X1 U2259 ( .A1(n793), .A2(n3828), .B1(n796), .B2(n3829), .ZN(n2193) );
  OAI221_X1 U2260 ( .B1(n40), .B2(n799), .C1(n264), .C2(n802), .A(n2194), .ZN(
        n2191) );
  AOI22_X1 U2261 ( .A1(n805), .A2(n1322), .B1(n808), .B2(n1355), .ZN(n2194) );
  OAI221_X1 U2262 ( .B1(n41), .B2(n811), .C1(n265), .C2(n814), .A(n2195), .ZN(
        n2190) );
  AOI22_X1 U2263 ( .A1(n817), .A2(n1183), .B1(n820), .B2(n1216), .ZN(n2195) );
  OAI221_X1 U2264 ( .B1(n42), .B2(n823), .C1(n266), .C2(n826), .A(n2196), .ZN(
        n2189) );
  AOI22_X1 U2265 ( .A1(n829), .A2(n1253), .B1(n832), .B2(n1286), .ZN(n2196) );
  NAND2_X1 U2266 ( .A1(n2197), .A2(n2198), .ZN(OUT1[3]) );
  NOR4_X1 U2267 ( .A1(n2199), .A2(n2200), .A3(n2201), .A4(n2202), .ZN(n2198)
         );
  OAI221_X1 U2268 ( .B1(n43), .B2(n739), .C1(n267), .C2(n742), .A(n2203), .ZN(
        n2202) );
  AOI22_X1 U2269 ( .A1(n745), .A2(n936), .B1(n748), .B2(n902), .ZN(n2203) );
  OAI221_X1 U2270 ( .B1(n44), .B2(n751), .C1(n268), .C2(n754), .A(n2204), .ZN(
        n2201) );
  AOI22_X1 U2271 ( .A1(n757), .A2(n1009), .B1(n760), .B2(n976), .ZN(n2204) );
  OAI221_X1 U2272 ( .B1(n45), .B2(n763), .C1(n269), .C2(n766), .A(n2205), .ZN(
        n2200) );
  AOI22_X1 U2273 ( .A1(n769), .A2(n1078), .B1(n772), .B2(n1045), .ZN(n2205) );
  OAI221_X1 U2274 ( .B1(n46), .B2(n775), .C1(n270), .C2(n778), .A(n2206), .ZN(
        n2199) );
  AOI22_X1 U2275 ( .A1(n781), .A2(n1147), .B1(n784), .B2(n1114), .ZN(n2206) );
  NOR4_X1 U2276 ( .A1(n2207), .A2(n2208), .A3(n2209), .A4(n2210), .ZN(n2197)
         );
  OAI221_X1 U2277 ( .B1(n3844), .B2(n787), .C1(n3845), .C2(n790), .A(n2211), 
        .ZN(n2210) );
  AOI22_X1 U2278 ( .A1(n793), .A2(n3846), .B1(n796), .B2(n3847), .ZN(n2211) );
  OAI221_X1 U2279 ( .B1(n47), .B2(n799), .C1(n271), .C2(n802), .A(n2212), .ZN(
        n2209) );
  AOI22_X1 U2280 ( .A1(n805), .A2(n1323), .B1(n808), .B2(n1356), .ZN(n2212) );
  OAI221_X1 U2281 ( .B1(n48), .B2(n811), .C1(n272), .C2(n814), .A(n2213), .ZN(
        n2208) );
  AOI22_X1 U2282 ( .A1(n817), .A2(n1184), .B1(n820), .B2(n1217), .ZN(n2213) );
  OAI221_X1 U2283 ( .B1(n49), .B2(n823), .C1(n273), .C2(n826), .A(n2214), .ZN(
        n2207) );
  AOI22_X1 U2284 ( .A1(n829), .A2(n1254), .B1(n832), .B2(n1287), .ZN(n2214) );
  NAND2_X1 U2285 ( .A1(n2215), .A2(n2216), .ZN(OUT1[31]) );
  NOR4_X1 U2286 ( .A1(n2217), .A2(n2218), .A3(n2219), .A4(n2220), .ZN(n2216)
         );
  OAI221_X1 U2287 ( .B1(n50), .B2(n739), .C1(n274), .C2(n742), .A(n2221), .ZN(
        n2220) );
  AOI22_X1 U2288 ( .A1(n745), .A2(n907), .B1(n748), .B2(n873), .ZN(n2221) );
  OAI221_X1 U2289 ( .B1(n51), .B2(n751), .C1(n275), .C2(n754), .A(n2222), .ZN(
        n2219) );
  AOI22_X1 U2290 ( .A1(n757), .A2(n980), .B1(n760), .B2(n947), .ZN(n2222) );
  OAI221_X1 U2291 ( .B1(n52), .B2(n763), .C1(n276), .C2(n766), .A(n2223), .ZN(
        n2218) );
  AOI22_X1 U2292 ( .A1(n769), .A2(n1049), .B1(n772), .B2(n1016), .ZN(n2223) );
  OAI221_X1 U2293 ( .B1(n53), .B2(n775), .C1(n277), .C2(n778), .A(n2224), .ZN(
        n2217) );
  AOI22_X1 U2294 ( .A1(n781), .A2(n1118), .B1(n784), .B2(n1085), .ZN(n2224) );
  NOR4_X1 U2295 ( .A1(n2225), .A2(n2226), .A3(n2227), .A4(n2228), .ZN(n2215)
         );
  OAI221_X1 U2296 ( .B1(n3862), .B2(n787), .C1(n3863), .C2(n790), .A(n2229), 
        .ZN(n2228) );
  AOI22_X1 U2297 ( .A1(n793), .A2(n3864), .B1(n796), .B2(n3865), .ZN(n2229) );
  OAI221_X1 U2298 ( .B1(n54), .B2(n799), .C1(n278), .C2(n802), .A(n2230), .ZN(
        n2227) );
  AOI22_X1 U2299 ( .A1(n805), .A2(n1294), .B1(n808), .B2(n1327), .ZN(n2230) );
  OAI221_X1 U2300 ( .B1(n55), .B2(n811), .C1(n279), .C2(n814), .A(n2231), .ZN(
        n2226) );
  AOI22_X1 U2301 ( .A1(n817), .A2(n1155), .B1(n820), .B2(n1188), .ZN(n2231) );
  OAI221_X1 U2302 ( .B1(n56), .B2(n823), .C1(n280), .C2(n826), .A(n2232), .ZN(
        n2225) );
  AOI22_X1 U2303 ( .A1(n829), .A2(n1225), .B1(n832), .B2(n1258), .ZN(n2232) );
  NAND2_X1 U2304 ( .A1(n2233), .A2(n2234), .ZN(OUT1[30]) );
  NOR4_X1 U2305 ( .A1(n2235), .A2(n2236), .A3(n2237), .A4(n2238), .ZN(n2234)
         );
  OAI221_X1 U2306 ( .B1(n57), .B2(n738), .C1(n281), .C2(n741), .A(n2239), .ZN(
        n2238) );
  AOI22_X1 U2307 ( .A1(n744), .A2(n909), .B1(n747), .B2(n875), .ZN(n2239) );
  OAI221_X1 U2308 ( .B1(n58), .B2(n750), .C1(n282), .C2(n753), .A(n2240), .ZN(
        n2237) );
  AOI22_X1 U2309 ( .A1(n756), .A2(n982), .B1(n759), .B2(n949), .ZN(n2240) );
  OAI221_X1 U2310 ( .B1(n59), .B2(n762), .C1(n283), .C2(n765), .A(n2241), .ZN(
        n2236) );
  AOI22_X1 U2311 ( .A1(n768), .A2(n1051), .B1(n771), .B2(n1018), .ZN(n2241) );
  OAI221_X1 U2312 ( .B1(n60), .B2(n774), .C1(n284), .C2(n777), .A(n2242), .ZN(
        n2235) );
  AOI22_X1 U2313 ( .A1(n780), .A2(n1120), .B1(n783), .B2(n1087), .ZN(n2242) );
  NOR4_X1 U2314 ( .A1(n2243), .A2(n2244), .A3(n2245), .A4(n2246), .ZN(n2233)
         );
  OAI221_X1 U2315 ( .B1(n3880), .B2(n786), .C1(n3881), .C2(n789), .A(n2247), 
        .ZN(n2246) );
  AOI22_X1 U2316 ( .A1(n792), .A2(n3882), .B1(n795), .B2(n3883), .ZN(n2247) );
  OAI221_X1 U2317 ( .B1(n61), .B2(n798), .C1(n285), .C2(n801), .A(n2248), .ZN(
        n2245) );
  AOI22_X1 U2318 ( .A1(n804), .A2(n1296), .B1(n807), .B2(n1329), .ZN(n2248) );
  OAI221_X1 U2319 ( .B1(n62), .B2(n810), .C1(n286), .C2(n813), .A(n2249), .ZN(
        n2244) );
  AOI22_X1 U2320 ( .A1(n816), .A2(n1157), .B1(n819), .B2(n1190), .ZN(n2249) );
  OAI221_X1 U2321 ( .B1(n63), .B2(n822), .C1(n287), .C2(n825), .A(n2250), .ZN(
        n2243) );
  AOI22_X1 U2322 ( .A1(n828), .A2(n1227), .B1(n831), .B2(n1260), .ZN(n2250) );
  NAND2_X1 U2323 ( .A1(n2251), .A2(n2252), .ZN(OUT1[2]) );
  NOR4_X1 U2324 ( .A1(n2253), .A2(n2254), .A3(n2255), .A4(n2256), .ZN(n2252)
         );
  OAI221_X1 U2325 ( .B1(n64), .B2(n738), .C1(n288), .C2(n741), .A(n2257), .ZN(
        n2256) );
  AOI22_X1 U2326 ( .A1(n744), .A2(n937), .B1(n747), .B2(n903), .ZN(n2257) );
  OAI221_X1 U2327 ( .B1(n65), .B2(n750), .C1(n289), .C2(n753), .A(n2258), .ZN(
        n2255) );
  AOI22_X1 U2328 ( .A1(n756), .A2(n1010), .B1(n759), .B2(n977), .ZN(n2258) );
  OAI221_X1 U2329 ( .B1(n66), .B2(n762), .C1(n290), .C2(n765), .A(n2259), .ZN(
        n2254) );
  AOI22_X1 U2330 ( .A1(n768), .A2(n1079), .B1(n771), .B2(n1046), .ZN(n2259) );
  OAI221_X1 U2331 ( .B1(n67), .B2(n774), .C1(n291), .C2(n777), .A(n2260), .ZN(
        n2253) );
  AOI22_X1 U2332 ( .A1(n780), .A2(n1148), .B1(n783), .B2(n1115), .ZN(n2260) );
  NOR4_X1 U2333 ( .A1(n2261), .A2(n2262), .A3(n2263), .A4(n2264), .ZN(n2251)
         );
  OAI221_X1 U2334 ( .B1(n3898), .B2(n786), .C1(n3899), .C2(n789), .A(n2265), 
        .ZN(n2264) );
  AOI22_X1 U2335 ( .A1(n792), .A2(n3900), .B1(n795), .B2(n3901), .ZN(n2265) );
  OAI221_X1 U2336 ( .B1(n68), .B2(n798), .C1(n292), .C2(n801), .A(n2266), .ZN(
        n2263) );
  AOI22_X1 U2337 ( .A1(n804), .A2(n1324), .B1(n807), .B2(n1357), .ZN(n2266) );
  OAI221_X1 U2338 ( .B1(n69), .B2(n810), .C1(n293), .C2(n813), .A(n2267), .ZN(
        n2262) );
  AOI22_X1 U2339 ( .A1(n816), .A2(n1185), .B1(n819), .B2(n1218), .ZN(n2267) );
  OAI221_X1 U2340 ( .B1(n70), .B2(n822), .C1(n294), .C2(n825), .A(n2268), .ZN(
        n2261) );
  AOI22_X1 U2341 ( .A1(n828), .A2(n1255), .B1(n831), .B2(n1288), .ZN(n2268) );
  NAND2_X1 U2342 ( .A1(n2269), .A2(n2270), .ZN(OUT1[29]) );
  NOR4_X1 U2343 ( .A1(n2271), .A2(n2272), .A3(n2273), .A4(n2274), .ZN(n2270)
         );
  OAI221_X1 U2344 ( .B1(n71), .B2(n738), .C1(n295), .C2(n741), .A(n2275), .ZN(
        n2274) );
  AOI22_X1 U2345 ( .A1(n744), .A2(n910), .B1(n747), .B2(n876), .ZN(n2275) );
  OAI221_X1 U2346 ( .B1(n72), .B2(n750), .C1(n296), .C2(n753), .A(n2276), .ZN(
        n2273) );
  AOI22_X1 U2347 ( .A1(n756), .A2(n983), .B1(n759), .B2(n950), .ZN(n2276) );
  OAI221_X1 U2348 ( .B1(n73), .B2(n762), .C1(n297), .C2(n765), .A(n2277), .ZN(
        n2272) );
  AOI22_X1 U2349 ( .A1(n768), .A2(n1052), .B1(n771), .B2(n1019), .ZN(n2277) );
  OAI221_X1 U2350 ( .B1(n74), .B2(n774), .C1(n298), .C2(n777), .A(n2278), .ZN(
        n2271) );
  AOI22_X1 U2351 ( .A1(n780), .A2(n1121), .B1(n783), .B2(n1088), .ZN(n2278) );
  NOR4_X1 U2352 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n2269)
         );
  OAI221_X1 U2353 ( .B1(n3916), .B2(n786), .C1(n3917), .C2(n789), .A(n2283), 
        .ZN(n2282) );
  AOI22_X1 U2354 ( .A1(n792), .A2(n3918), .B1(n795), .B2(n3919), .ZN(n2283) );
  OAI221_X1 U2355 ( .B1(n75), .B2(n798), .C1(n299), .C2(n801), .A(n2284), .ZN(
        n2281) );
  AOI22_X1 U2356 ( .A1(n804), .A2(n1297), .B1(n807), .B2(n1330), .ZN(n2284) );
  OAI221_X1 U2357 ( .B1(n76), .B2(n810), .C1(n300), .C2(n813), .A(n2285), .ZN(
        n2280) );
  AOI22_X1 U2358 ( .A1(n816), .A2(n1158), .B1(n819), .B2(n1191), .ZN(n2285) );
  OAI221_X1 U2359 ( .B1(n77), .B2(n822), .C1(n301), .C2(n825), .A(n2286), .ZN(
        n2279) );
  AOI22_X1 U2360 ( .A1(n828), .A2(n1228), .B1(n831), .B2(n1261), .ZN(n2286) );
  NAND2_X1 U2361 ( .A1(n2287), .A2(n2288), .ZN(OUT1[28]) );
  NOR4_X1 U2362 ( .A1(n2289), .A2(n2290), .A3(n2291), .A4(n2292), .ZN(n2288)
         );
  OAI221_X1 U2363 ( .B1(n78), .B2(n738), .C1(n302), .C2(n741), .A(n2293), .ZN(
        n2292) );
  AOI22_X1 U2364 ( .A1(n744), .A2(n911), .B1(n747), .B2(n877), .ZN(n2293) );
  OAI221_X1 U2365 ( .B1(n79), .B2(n750), .C1(n303), .C2(n753), .A(n2294), .ZN(
        n2291) );
  AOI22_X1 U2366 ( .A1(n756), .A2(n984), .B1(n759), .B2(n951), .ZN(n2294) );
  OAI221_X1 U2367 ( .B1(n80), .B2(n762), .C1(n304), .C2(n765), .A(n2295), .ZN(
        n2290) );
  AOI22_X1 U2368 ( .A1(n768), .A2(n1053), .B1(n771), .B2(n1020), .ZN(n2295) );
  OAI221_X1 U2369 ( .B1(n81), .B2(n774), .C1(n305), .C2(n777), .A(n2296), .ZN(
        n2289) );
  AOI22_X1 U2370 ( .A1(n780), .A2(n1122), .B1(n783), .B2(n1089), .ZN(n2296) );
  NOR4_X1 U2371 ( .A1(n2297), .A2(n2298), .A3(n2299), .A4(n2300), .ZN(n2287)
         );
  OAI221_X1 U2372 ( .B1(n3934), .B2(n786), .C1(n3935), .C2(n789), .A(n2301), 
        .ZN(n2300) );
  AOI22_X1 U2373 ( .A1(n792), .A2(n3936), .B1(n795), .B2(n3937), .ZN(n2301) );
  OAI221_X1 U2374 ( .B1(n82), .B2(n798), .C1(n306), .C2(n801), .A(n2302), .ZN(
        n2299) );
  AOI22_X1 U2375 ( .A1(n804), .A2(n1298), .B1(n807), .B2(n1331), .ZN(n2302) );
  OAI221_X1 U2376 ( .B1(n83), .B2(n810), .C1(n307), .C2(n813), .A(n2303), .ZN(
        n2298) );
  AOI22_X1 U2377 ( .A1(n816), .A2(n1159), .B1(n819), .B2(n1192), .ZN(n2303) );
  OAI221_X1 U2378 ( .B1(n84), .B2(n822), .C1(n308), .C2(n825), .A(n2304), .ZN(
        n2297) );
  AOI22_X1 U2379 ( .A1(n828), .A2(n1229), .B1(n831), .B2(n1262), .ZN(n2304) );
  NAND2_X1 U2380 ( .A1(n2305), .A2(n2306), .ZN(OUT1[27]) );
  NOR4_X1 U2381 ( .A1(n2307), .A2(n2308), .A3(n2309), .A4(n2310), .ZN(n2306)
         );
  OAI221_X1 U2382 ( .B1(n85), .B2(n738), .C1(n309), .C2(n741), .A(n2311), .ZN(
        n2310) );
  AOI22_X1 U2383 ( .A1(n744), .A2(n912), .B1(n747), .B2(n878), .ZN(n2311) );
  OAI221_X1 U2384 ( .B1(n86), .B2(n750), .C1(n310), .C2(n753), .A(n2312), .ZN(
        n2309) );
  AOI22_X1 U2385 ( .A1(n756), .A2(n985), .B1(n759), .B2(n952), .ZN(n2312) );
  OAI221_X1 U2386 ( .B1(n87), .B2(n762), .C1(n311), .C2(n765), .A(n2313), .ZN(
        n2308) );
  AOI22_X1 U2387 ( .A1(n768), .A2(n1054), .B1(n771), .B2(n1021), .ZN(n2313) );
  OAI221_X1 U2388 ( .B1(n88), .B2(n774), .C1(n312), .C2(n777), .A(n2314), .ZN(
        n2307) );
  AOI22_X1 U2389 ( .A1(n780), .A2(n1123), .B1(n783), .B2(n1090), .ZN(n2314) );
  NOR4_X1 U2390 ( .A1(n2315), .A2(n2316), .A3(n2317), .A4(n2318), .ZN(n2305)
         );
  OAI221_X1 U2391 ( .B1(n3952), .B2(n786), .C1(n3953), .C2(n789), .A(n2319), 
        .ZN(n2318) );
  AOI22_X1 U2392 ( .A1(n792), .A2(n3954), .B1(n795), .B2(n3955), .ZN(n2319) );
  OAI221_X1 U2393 ( .B1(n89), .B2(n798), .C1(n313), .C2(n801), .A(n2320), .ZN(
        n2317) );
  AOI22_X1 U2394 ( .A1(n804), .A2(n1299), .B1(n807), .B2(n1332), .ZN(n2320) );
  OAI221_X1 U2395 ( .B1(n90), .B2(n810), .C1(n314), .C2(n813), .A(n2321), .ZN(
        n2316) );
  AOI22_X1 U2396 ( .A1(n816), .A2(n1160), .B1(n819), .B2(n1193), .ZN(n2321) );
  OAI221_X1 U2397 ( .B1(n91), .B2(n822), .C1(n315), .C2(n825), .A(n2322), .ZN(
        n2315) );
  AOI22_X1 U2398 ( .A1(n828), .A2(n1230), .B1(n831), .B2(n1263), .ZN(n2322) );
  NAND2_X1 U2399 ( .A1(n2323), .A2(n2324), .ZN(OUT1[26]) );
  NOR4_X1 U2400 ( .A1(n2325), .A2(n2326), .A3(n2327), .A4(n2328), .ZN(n2324)
         );
  OAI221_X1 U2401 ( .B1(n92), .B2(n738), .C1(n316), .C2(n741), .A(n2329), .ZN(
        n2328) );
  AOI22_X1 U2402 ( .A1(n744), .A2(n913), .B1(n747), .B2(n879), .ZN(n2329) );
  OAI221_X1 U2403 ( .B1(n93), .B2(n750), .C1(n317), .C2(n753), .A(n2330), .ZN(
        n2327) );
  AOI22_X1 U2404 ( .A1(n756), .A2(n986), .B1(n759), .B2(n953), .ZN(n2330) );
  OAI221_X1 U2405 ( .B1(n94), .B2(n762), .C1(n318), .C2(n765), .A(n2331), .ZN(
        n2326) );
  AOI22_X1 U2406 ( .A1(n768), .A2(n1055), .B1(n771), .B2(n1022), .ZN(n2331) );
  OAI221_X1 U2407 ( .B1(n95), .B2(n774), .C1(n319), .C2(n777), .A(n2332), .ZN(
        n2325) );
  AOI22_X1 U2408 ( .A1(n780), .A2(n1124), .B1(n783), .B2(n1091), .ZN(n2332) );
  NOR4_X1 U2409 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(n2323)
         );
  OAI221_X1 U2410 ( .B1(n3970), .B2(n786), .C1(n3971), .C2(n789), .A(n2337), 
        .ZN(n2336) );
  AOI22_X1 U2411 ( .A1(n792), .A2(n3972), .B1(n795), .B2(n3973), .ZN(n2337) );
  OAI221_X1 U2412 ( .B1(n96), .B2(n798), .C1(n320), .C2(n801), .A(n2338), .ZN(
        n2335) );
  AOI22_X1 U2413 ( .A1(n804), .A2(n1300), .B1(n807), .B2(n1333), .ZN(n2338) );
  OAI221_X1 U2414 ( .B1(n97), .B2(n810), .C1(n321), .C2(n813), .A(n2339), .ZN(
        n2334) );
  AOI22_X1 U2415 ( .A1(n816), .A2(n1161), .B1(n819), .B2(n1194), .ZN(n2339) );
  OAI221_X1 U2416 ( .B1(n98), .B2(n822), .C1(n322), .C2(n825), .A(n2340), .ZN(
        n2333) );
  AOI22_X1 U2417 ( .A1(n828), .A2(n1231), .B1(n831), .B2(n1264), .ZN(n2340) );
  NAND2_X1 U2418 ( .A1(n2341), .A2(n2342), .ZN(OUT1[25]) );
  NOR4_X1 U2419 ( .A1(n2343), .A2(n2344), .A3(n2345), .A4(n2346), .ZN(n2342)
         );
  OAI221_X1 U2420 ( .B1(n99), .B2(n738), .C1(n323), .C2(n741), .A(n2347), .ZN(
        n2346) );
  AOI22_X1 U2421 ( .A1(n744), .A2(n914), .B1(n747), .B2(n880), .ZN(n2347) );
  OAI221_X1 U2422 ( .B1(n100), .B2(n750), .C1(n324), .C2(n753), .A(n2348), 
        .ZN(n2345) );
  AOI22_X1 U2423 ( .A1(n756), .A2(n987), .B1(n759), .B2(n954), .ZN(n2348) );
  OAI221_X1 U2424 ( .B1(n101), .B2(n762), .C1(n325), .C2(n765), .A(n2349), 
        .ZN(n2344) );
  AOI22_X1 U2425 ( .A1(n768), .A2(n1056), .B1(n771), .B2(n1023), .ZN(n2349) );
  OAI221_X1 U2426 ( .B1(n102), .B2(n774), .C1(n326), .C2(n777), .A(n2350), 
        .ZN(n2343) );
  AOI22_X1 U2427 ( .A1(n780), .A2(n1125), .B1(n783), .B2(n1092), .ZN(n2350) );
  NOR4_X1 U2428 ( .A1(n2351), .A2(n2352), .A3(n2353), .A4(n2354), .ZN(n2341)
         );
  OAI221_X1 U2429 ( .B1(n3988), .B2(n786), .C1(n3989), .C2(n789), .A(n2355), 
        .ZN(n2354) );
  AOI22_X1 U2430 ( .A1(n792), .A2(n3990), .B1(n795), .B2(n3991), .ZN(n2355) );
  OAI221_X1 U2431 ( .B1(n103), .B2(n798), .C1(n327), .C2(n801), .A(n2356), 
        .ZN(n2353) );
  AOI22_X1 U2432 ( .A1(n804), .A2(n1301), .B1(n807), .B2(n1334), .ZN(n2356) );
  OAI221_X1 U2433 ( .B1(n104), .B2(n810), .C1(n328), .C2(n813), .A(n2357), 
        .ZN(n2352) );
  AOI22_X1 U2434 ( .A1(n816), .A2(n1162), .B1(n819), .B2(n1195), .ZN(n2357) );
  OAI221_X1 U2435 ( .B1(n105), .B2(n822), .C1(n329), .C2(n825), .A(n2358), 
        .ZN(n2351) );
  AOI22_X1 U2436 ( .A1(n828), .A2(n1232), .B1(n831), .B2(n1265), .ZN(n2358) );
  NAND2_X1 U2437 ( .A1(n2359), .A2(n2360), .ZN(OUT1[24]) );
  NOR4_X1 U2438 ( .A1(n2361), .A2(n2362), .A3(n2363), .A4(n2364), .ZN(n2360)
         );
  OAI221_X1 U2439 ( .B1(n106), .B2(n738), .C1(n330), .C2(n741), .A(n2365), 
        .ZN(n2364) );
  AOI22_X1 U2440 ( .A1(n744), .A2(n915), .B1(n747), .B2(n881), .ZN(n2365) );
  OAI221_X1 U2441 ( .B1(n107), .B2(n750), .C1(n331), .C2(n753), .A(n2366), 
        .ZN(n2363) );
  AOI22_X1 U2442 ( .A1(n756), .A2(n988), .B1(n759), .B2(n955), .ZN(n2366) );
  OAI221_X1 U2443 ( .B1(n108), .B2(n762), .C1(n332), .C2(n765), .A(n2367), 
        .ZN(n2362) );
  AOI22_X1 U2444 ( .A1(n768), .A2(n1057), .B1(n771), .B2(n1024), .ZN(n2367) );
  OAI221_X1 U2445 ( .B1(n109), .B2(n774), .C1(n333), .C2(n777), .A(n2368), 
        .ZN(n2361) );
  AOI22_X1 U2446 ( .A1(n780), .A2(n1126), .B1(n783), .B2(n1093), .ZN(n2368) );
  NOR4_X1 U2447 ( .A1(n2369), .A2(n2370), .A3(n2371), .A4(n2372), .ZN(n2359)
         );
  OAI221_X1 U2448 ( .B1(n4006), .B2(n786), .C1(n4007), .C2(n789), .A(n2373), 
        .ZN(n2372) );
  AOI22_X1 U2449 ( .A1(n792), .A2(n4008), .B1(n795), .B2(n4009), .ZN(n2373) );
  OAI221_X1 U2450 ( .B1(n110), .B2(n798), .C1(n334), .C2(n801), .A(n2374), 
        .ZN(n2371) );
  AOI22_X1 U2451 ( .A1(n804), .A2(n1302), .B1(n807), .B2(n1335), .ZN(n2374) );
  OAI221_X1 U2452 ( .B1(n111), .B2(n810), .C1(n335), .C2(n813), .A(n2375), 
        .ZN(n2370) );
  AOI22_X1 U2453 ( .A1(n816), .A2(n1163), .B1(n819), .B2(n1196), .ZN(n2375) );
  OAI221_X1 U2454 ( .B1(n112), .B2(n822), .C1(n336), .C2(n825), .A(n2376), 
        .ZN(n2369) );
  AOI22_X1 U2455 ( .A1(n828), .A2(n1233), .B1(n831), .B2(n1266), .ZN(n2376) );
  NAND2_X1 U2456 ( .A1(n2377), .A2(n2378), .ZN(OUT1[23]) );
  NOR4_X1 U2457 ( .A1(n2379), .A2(n2380), .A3(n2381), .A4(n2382), .ZN(n2378)
         );
  OAI221_X1 U2458 ( .B1(n113), .B2(n738), .C1(n337), .C2(n741), .A(n2383), 
        .ZN(n2382) );
  AOI22_X1 U2459 ( .A1(n744), .A2(n916), .B1(n747), .B2(n882), .ZN(n2383) );
  OAI221_X1 U2460 ( .B1(n114), .B2(n750), .C1(n338), .C2(n753), .A(n2384), 
        .ZN(n2381) );
  AOI22_X1 U2461 ( .A1(n756), .A2(n989), .B1(n759), .B2(n956), .ZN(n2384) );
  OAI221_X1 U2462 ( .B1(n115), .B2(n762), .C1(n339), .C2(n765), .A(n2385), 
        .ZN(n2380) );
  AOI22_X1 U2463 ( .A1(n768), .A2(n1058), .B1(n771), .B2(n1025), .ZN(n2385) );
  OAI221_X1 U2464 ( .B1(n116), .B2(n774), .C1(n340), .C2(n777), .A(n2386), 
        .ZN(n2379) );
  AOI22_X1 U2465 ( .A1(n780), .A2(n1127), .B1(n783), .B2(n1094), .ZN(n2386) );
  NOR4_X1 U2466 ( .A1(n2387), .A2(n2388), .A3(n2389), .A4(n2390), .ZN(n2377)
         );
  OAI221_X1 U2467 ( .B1(n4024), .B2(n786), .C1(n4025), .C2(n789), .A(n2391), 
        .ZN(n2390) );
  AOI22_X1 U2468 ( .A1(n792), .A2(n4026), .B1(n795), .B2(n4027), .ZN(n2391) );
  OAI221_X1 U2469 ( .B1(n117), .B2(n798), .C1(n341), .C2(n801), .A(n2392), 
        .ZN(n2389) );
  AOI22_X1 U2470 ( .A1(n804), .A2(n1303), .B1(n807), .B2(n1336), .ZN(n2392) );
  OAI221_X1 U2471 ( .B1(n118), .B2(n810), .C1(n342), .C2(n813), .A(n2393), 
        .ZN(n2388) );
  AOI22_X1 U2472 ( .A1(n816), .A2(n1164), .B1(n819), .B2(n1197), .ZN(n2393) );
  OAI221_X1 U2473 ( .B1(n119), .B2(n822), .C1(n343), .C2(n825), .A(n2394), 
        .ZN(n2387) );
  AOI22_X1 U2474 ( .A1(n828), .A2(n1234), .B1(n831), .B2(n1267), .ZN(n2394) );
  NAND2_X1 U2475 ( .A1(n2395), .A2(n2396), .ZN(OUT1[22]) );
  NOR4_X1 U2476 ( .A1(n2397), .A2(n2398), .A3(n2399), .A4(n2400), .ZN(n2396)
         );
  OAI221_X1 U2477 ( .B1(n120), .B2(n738), .C1(n344), .C2(n741), .A(n2401), 
        .ZN(n2400) );
  AOI22_X1 U2478 ( .A1(n744), .A2(n917), .B1(n747), .B2(n883), .ZN(n2401) );
  OAI221_X1 U2479 ( .B1(n121), .B2(n750), .C1(n345), .C2(n753), .A(n2402), 
        .ZN(n2399) );
  AOI22_X1 U2480 ( .A1(n756), .A2(n990), .B1(n759), .B2(n957), .ZN(n2402) );
  OAI221_X1 U2481 ( .B1(n122), .B2(n762), .C1(n346), .C2(n765), .A(n2403), 
        .ZN(n2398) );
  AOI22_X1 U2482 ( .A1(n768), .A2(n1059), .B1(n771), .B2(n1026), .ZN(n2403) );
  OAI221_X1 U2483 ( .B1(n123), .B2(n774), .C1(n347), .C2(n777), .A(n2404), 
        .ZN(n2397) );
  AOI22_X1 U2484 ( .A1(n780), .A2(n1128), .B1(n783), .B2(n1095), .ZN(n2404) );
  NOR4_X1 U2485 ( .A1(n2405), .A2(n2406), .A3(n2407), .A4(n2408), .ZN(n2395)
         );
  OAI221_X1 U2486 ( .B1(n4042), .B2(n786), .C1(n4043), .C2(n789), .A(n2409), 
        .ZN(n2408) );
  AOI22_X1 U2487 ( .A1(n792), .A2(n4044), .B1(n795), .B2(n4045), .ZN(n2409) );
  OAI221_X1 U2488 ( .B1(n124), .B2(n798), .C1(n348), .C2(n801), .A(n2410), 
        .ZN(n2407) );
  AOI22_X1 U2489 ( .A1(n804), .A2(n1304), .B1(n807), .B2(n1337), .ZN(n2410) );
  OAI221_X1 U2490 ( .B1(n125), .B2(n810), .C1(n349), .C2(n813), .A(n2411), 
        .ZN(n2406) );
  AOI22_X1 U2491 ( .A1(n816), .A2(n1165), .B1(n819), .B2(n1198), .ZN(n2411) );
  OAI221_X1 U2492 ( .B1(n126), .B2(n822), .C1(n350), .C2(n825), .A(n2412), 
        .ZN(n2405) );
  AOI22_X1 U2493 ( .A1(n828), .A2(n1235), .B1(n831), .B2(n1268), .ZN(n2412) );
  NAND2_X1 U2494 ( .A1(n2413), .A2(n2414), .ZN(OUT1[21]) );
  NOR4_X1 U2495 ( .A1(n2415), .A2(n2416), .A3(n2417), .A4(n2418), .ZN(n2414)
         );
  OAI221_X1 U2496 ( .B1(n127), .B2(n738), .C1(n351), .C2(n741), .A(n2419), 
        .ZN(n2418) );
  AOI22_X1 U2497 ( .A1(n744), .A2(n918), .B1(n747), .B2(n884), .ZN(n2419) );
  OAI221_X1 U2498 ( .B1(n128), .B2(n750), .C1(n352), .C2(n753), .A(n2420), 
        .ZN(n2417) );
  AOI22_X1 U2499 ( .A1(n756), .A2(n991), .B1(n759), .B2(n958), .ZN(n2420) );
  OAI221_X1 U2500 ( .B1(n129), .B2(n762), .C1(n353), .C2(n765), .A(n2421), 
        .ZN(n2416) );
  AOI22_X1 U2501 ( .A1(n768), .A2(n1060), .B1(n771), .B2(n1027), .ZN(n2421) );
  OAI221_X1 U2502 ( .B1(n130), .B2(n774), .C1(n354), .C2(n777), .A(n2422), 
        .ZN(n2415) );
  AOI22_X1 U2503 ( .A1(n780), .A2(n1129), .B1(n783), .B2(n1096), .ZN(n2422) );
  NOR4_X1 U2504 ( .A1(n2423), .A2(n2424), .A3(n2425), .A4(n2426), .ZN(n2413)
         );
  OAI221_X1 U2505 ( .B1(n4060), .B2(n786), .C1(n4061), .C2(n789), .A(n2427), 
        .ZN(n2426) );
  AOI22_X1 U2506 ( .A1(n792), .A2(n4062), .B1(n795), .B2(n4063), .ZN(n2427) );
  OAI221_X1 U2507 ( .B1(n131), .B2(n798), .C1(n355), .C2(n801), .A(n2428), 
        .ZN(n2425) );
  AOI22_X1 U2508 ( .A1(n804), .A2(n1305), .B1(n807), .B2(n1338), .ZN(n2428) );
  OAI221_X1 U2509 ( .B1(n132), .B2(n810), .C1(n356), .C2(n813), .A(n2429), 
        .ZN(n2424) );
  AOI22_X1 U2510 ( .A1(n816), .A2(n1166), .B1(n819), .B2(n1199), .ZN(n2429) );
  OAI221_X1 U2511 ( .B1(n133), .B2(n822), .C1(n357), .C2(n825), .A(n2430), 
        .ZN(n2423) );
  AOI22_X1 U2512 ( .A1(n828), .A2(n1236), .B1(n831), .B2(n1269), .ZN(n2430) );
  NAND2_X1 U2513 ( .A1(n2431), .A2(n2432), .ZN(OUT1[20]) );
  NOR4_X1 U2514 ( .A1(n2433), .A2(n2434), .A3(n2435), .A4(n2436), .ZN(n2432)
         );
  OAI221_X1 U2515 ( .B1(n134), .B2(n738), .C1(n358), .C2(n741), .A(n2437), 
        .ZN(n2436) );
  AOI22_X1 U2516 ( .A1(n744), .A2(n919), .B1(n747), .B2(n885), .ZN(n2437) );
  OAI221_X1 U2517 ( .B1(n135), .B2(n750), .C1(n359), .C2(n753), .A(n2438), 
        .ZN(n2435) );
  AOI22_X1 U2518 ( .A1(n756), .A2(n992), .B1(n759), .B2(n959), .ZN(n2438) );
  OAI221_X1 U2519 ( .B1(n136), .B2(n762), .C1(n360), .C2(n765), .A(n2439), 
        .ZN(n2434) );
  AOI22_X1 U2520 ( .A1(n768), .A2(n1061), .B1(n771), .B2(n1028), .ZN(n2439) );
  OAI221_X1 U2521 ( .B1(n137), .B2(n774), .C1(n361), .C2(n777), .A(n2440), 
        .ZN(n2433) );
  AOI22_X1 U2522 ( .A1(n780), .A2(n1130), .B1(n783), .B2(n1097), .ZN(n2440) );
  NOR4_X1 U2523 ( .A1(n2441), .A2(n2442), .A3(n2443), .A4(n2444), .ZN(n2431)
         );
  OAI221_X1 U2524 ( .B1(n4078), .B2(n786), .C1(n4079), .C2(n789), .A(n2445), 
        .ZN(n2444) );
  AOI22_X1 U2525 ( .A1(n792), .A2(n4080), .B1(n795), .B2(n4081), .ZN(n2445) );
  OAI221_X1 U2526 ( .B1(n138), .B2(n798), .C1(n362), .C2(n801), .A(n2446), 
        .ZN(n2443) );
  AOI22_X1 U2527 ( .A1(n804), .A2(n1306), .B1(n807), .B2(n1339), .ZN(n2446) );
  OAI221_X1 U2528 ( .B1(n139), .B2(n810), .C1(n363), .C2(n813), .A(n2447), 
        .ZN(n2442) );
  AOI22_X1 U2529 ( .A1(n816), .A2(n1167), .B1(n819), .B2(n1200), .ZN(n2447) );
  OAI221_X1 U2530 ( .B1(n140), .B2(n822), .C1(n364), .C2(n825), .A(n2448), 
        .ZN(n2441) );
  AOI22_X1 U2531 ( .A1(n828), .A2(n1237), .B1(n831), .B2(n1270), .ZN(n2448) );
  NAND2_X1 U2532 ( .A1(n2449), .A2(n2450), .ZN(OUT1[1]) );
  NOR4_X1 U2533 ( .A1(n2451), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(n2450)
         );
  OAI221_X1 U2534 ( .B1(n141), .B2(n737), .C1(n365), .C2(n740), .A(n2455), 
        .ZN(n2454) );
  AOI22_X1 U2535 ( .A1(n743), .A2(n938), .B1(n746), .B2(n904), .ZN(n2455) );
  OAI221_X1 U2536 ( .B1(n142), .B2(n749), .C1(n366), .C2(n752), .A(n2456), 
        .ZN(n2453) );
  AOI22_X1 U2537 ( .A1(n755), .A2(n1011), .B1(n758), .B2(n978), .ZN(n2456) );
  OAI221_X1 U2538 ( .B1(n143), .B2(n761), .C1(n367), .C2(n764), .A(n2457), 
        .ZN(n2452) );
  AOI22_X1 U2539 ( .A1(n767), .A2(n1080), .B1(n770), .B2(n1047), .ZN(n2457) );
  OAI221_X1 U2540 ( .B1(n144), .B2(n773), .C1(n368), .C2(n776), .A(n2458), 
        .ZN(n2451) );
  AOI22_X1 U2541 ( .A1(n779), .A2(n1149), .B1(n782), .B2(n1116), .ZN(n2458) );
  NOR4_X1 U2542 ( .A1(n2459), .A2(n2460), .A3(n2461), .A4(n2462), .ZN(n2449)
         );
  OAI221_X1 U2543 ( .B1(n4096), .B2(n785), .C1(n4097), .C2(n788), .A(n2463), 
        .ZN(n2462) );
  AOI22_X1 U2544 ( .A1(n791), .A2(n4098), .B1(n794), .B2(n4099), .ZN(n2463) );
  OAI221_X1 U2545 ( .B1(n145), .B2(n797), .C1(n369), .C2(n800), .A(n2464), 
        .ZN(n2461) );
  AOI22_X1 U2546 ( .A1(n803), .A2(n1325), .B1(n806), .B2(n1358), .ZN(n2464) );
  OAI221_X1 U2547 ( .B1(n146), .B2(n809), .C1(n370), .C2(n812), .A(n2465), 
        .ZN(n2460) );
  AOI22_X1 U2548 ( .A1(n815), .A2(n1186), .B1(n818), .B2(n1219), .ZN(n2465) );
  OAI221_X1 U2549 ( .B1(n147), .B2(n821), .C1(n371), .C2(n824), .A(n2466), 
        .ZN(n2459) );
  AOI22_X1 U2550 ( .A1(n827), .A2(n1256), .B1(n830), .B2(n1289), .ZN(n2466) );
  NAND2_X1 U2551 ( .A1(n2467), .A2(n2468), .ZN(OUT1[19]) );
  NOR4_X1 U2552 ( .A1(n2469), .A2(n2470), .A3(n2471), .A4(n2472), .ZN(n2468)
         );
  OAI221_X1 U2553 ( .B1(n148), .B2(n737), .C1(n372), .C2(n740), .A(n2473), 
        .ZN(n2472) );
  AOI22_X1 U2554 ( .A1(n743), .A2(n920), .B1(n746), .B2(n886), .ZN(n2473) );
  OAI221_X1 U2555 ( .B1(n149), .B2(n749), .C1(n373), .C2(n752), .A(n2474), 
        .ZN(n2471) );
  AOI22_X1 U2556 ( .A1(n755), .A2(n993), .B1(n758), .B2(n960), .ZN(n2474) );
  OAI221_X1 U2557 ( .B1(n150), .B2(n761), .C1(n374), .C2(n764), .A(n2475), 
        .ZN(n2470) );
  AOI22_X1 U2558 ( .A1(n767), .A2(n1062), .B1(n770), .B2(n1029), .ZN(n2475) );
  OAI221_X1 U2559 ( .B1(n151), .B2(n773), .C1(n375), .C2(n776), .A(n2476), 
        .ZN(n2469) );
  AOI22_X1 U2560 ( .A1(n779), .A2(n1131), .B1(n782), .B2(n1098), .ZN(n2476) );
  NOR4_X1 U2561 ( .A1(n2477), .A2(n2478), .A3(n2479), .A4(n2480), .ZN(n2467)
         );
  OAI221_X1 U2562 ( .B1(n4114), .B2(n785), .C1(n4115), .C2(n788), .A(n2481), 
        .ZN(n2480) );
  AOI22_X1 U2563 ( .A1(n791), .A2(n4116), .B1(n794), .B2(n4117), .ZN(n2481) );
  OAI221_X1 U2564 ( .B1(n152), .B2(n797), .C1(n376), .C2(n800), .A(n2482), 
        .ZN(n2479) );
  AOI22_X1 U2565 ( .A1(n803), .A2(n1307), .B1(n806), .B2(n1340), .ZN(n2482) );
  OAI221_X1 U2566 ( .B1(n153), .B2(n809), .C1(n377), .C2(n812), .A(n2483), 
        .ZN(n2478) );
  AOI22_X1 U2567 ( .A1(n815), .A2(n1168), .B1(n818), .B2(n1201), .ZN(n2483) );
  OAI221_X1 U2568 ( .B1(n154), .B2(n821), .C1(n378), .C2(n824), .A(n2484), 
        .ZN(n2477) );
  AOI22_X1 U2569 ( .A1(n827), .A2(n1238), .B1(n830), .B2(n1271), .ZN(n2484) );
  NAND2_X1 U2570 ( .A1(n2485), .A2(n2486), .ZN(OUT1[18]) );
  NOR4_X1 U2571 ( .A1(n2487), .A2(n2488), .A3(n2489), .A4(n2490), .ZN(n2486)
         );
  OAI221_X1 U2572 ( .B1(n155), .B2(n737), .C1(n379), .C2(n740), .A(n2491), 
        .ZN(n2490) );
  AOI22_X1 U2573 ( .A1(n743), .A2(n921), .B1(n746), .B2(n887), .ZN(n2491) );
  OAI221_X1 U2574 ( .B1(n156), .B2(n749), .C1(n380), .C2(n752), .A(n2492), 
        .ZN(n2489) );
  AOI22_X1 U2575 ( .A1(n755), .A2(n994), .B1(n758), .B2(n961), .ZN(n2492) );
  OAI221_X1 U2576 ( .B1(n157), .B2(n761), .C1(n381), .C2(n764), .A(n2493), 
        .ZN(n2488) );
  AOI22_X1 U2577 ( .A1(n767), .A2(n1063), .B1(n770), .B2(n1030), .ZN(n2493) );
  OAI221_X1 U2578 ( .B1(n158), .B2(n773), .C1(n382), .C2(n776), .A(n2494), 
        .ZN(n2487) );
  AOI22_X1 U2579 ( .A1(n779), .A2(n1132), .B1(n782), .B2(n1099), .ZN(n2494) );
  NOR4_X1 U2580 ( .A1(n2495), .A2(n2496), .A3(n2497), .A4(n2498), .ZN(n2485)
         );
  OAI221_X1 U2581 ( .B1(n4132), .B2(n785), .C1(n4133), .C2(n788), .A(n2499), 
        .ZN(n2498) );
  AOI22_X1 U2582 ( .A1(n791), .A2(n4134), .B1(n794), .B2(n4135), .ZN(n2499) );
  OAI221_X1 U2583 ( .B1(n159), .B2(n797), .C1(n383), .C2(n800), .A(n2500), 
        .ZN(n2497) );
  AOI22_X1 U2584 ( .A1(n803), .A2(n1308), .B1(n806), .B2(n1341), .ZN(n2500) );
  OAI221_X1 U2585 ( .B1(n160), .B2(n809), .C1(n384), .C2(n812), .A(n2501), 
        .ZN(n2496) );
  AOI22_X1 U2586 ( .A1(n815), .A2(n1169), .B1(n818), .B2(n1202), .ZN(n2501) );
  OAI221_X1 U2587 ( .B1(n161), .B2(n821), .C1(n385), .C2(n824), .A(n2502), 
        .ZN(n2495) );
  AOI22_X1 U2588 ( .A1(n827), .A2(n1239), .B1(n830), .B2(n1272), .ZN(n2502) );
  NAND2_X1 U2589 ( .A1(n2503), .A2(n2504), .ZN(OUT1[17]) );
  NOR4_X1 U2590 ( .A1(n2505), .A2(n2506), .A3(n2507), .A4(n2508), .ZN(n2504)
         );
  OAI221_X1 U2591 ( .B1(n162), .B2(n737), .C1(n386), .C2(n740), .A(n2509), 
        .ZN(n2508) );
  AOI22_X1 U2592 ( .A1(n743), .A2(n922), .B1(n746), .B2(n888), .ZN(n2509) );
  OAI221_X1 U2593 ( .B1(n163), .B2(n749), .C1(n387), .C2(n752), .A(n2510), 
        .ZN(n2507) );
  AOI22_X1 U2594 ( .A1(n755), .A2(n995), .B1(n758), .B2(n962), .ZN(n2510) );
  OAI221_X1 U2595 ( .B1(n164), .B2(n761), .C1(n388), .C2(n764), .A(n2511), 
        .ZN(n2506) );
  AOI22_X1 U2596 ( .A1(n767), .A2(n1064), .B1(n770), .B2(n1031), .ZN(n2511) );
  OAI221_X1 U2597 ( .B1(n165), .B2(n773), .C1(n389), .C2(n776), .A(n2512), 
        .ZN(n2505) );
  AOI22_X1 U2598 ( .A1(n779), .A2(n1133), .B1(n782), .B2(n1100), .ZN(n2512) );
  NOR4_X1 U2599 ( .A1(n2513), .A2(n2514), .A3(n2515), .A4(n2516), .ZN(n2503)
         );
  OAI221_X1 U2600 ( .B1(n4150), .B2(n785), .C1(n4151), .C2(n788), .A(n2517), 
        .ZN(n2516) );
  AOI22_X1 U2601 ( .A1(n791), .A2(n4152), .B1(n794), .B2(n4153), .ZN(n2517) );
  OAI221_X1 U2602 ( .B1(n166), .B2(n797), .C1(n390), .C2(n800), .A(n2518), 
        .ZN(n2515) );
  AOI22_X1 U2603 ( .A1(n803), .A2(n1309), .B1(n806), .B2(n1342), .ZN(n2518) );
  OAI221_X1 U2604 ( .B1(n167), .B2(n809), .C1(n391), .C2(n812), .A(n2519), 
        .ZN(n2514) );
  AOI22_X1 U2605 ( .A1(n815), .A2(n1170), .B1(n818), .B2(n1203), .ZN(n2519) );
  OAI221_X1 U2606 ( .B1(n168), .B2(n821), .C1(n392), .C2(n824), .A(n2520), 
        .ZN(n2513) );
  AOI22_X1 U2607 ( .A1(n827), .A2(n1240), .B1(n830), .B2(n1273), .ZN(n2520) );
  NAND2_X1 U2608 ( .A1(n2521), .A2(n2522), .ZN(OUT1[16]) );
  NOR4_X1 U2609 ( .A1(n2523), .A2(n2524), .A3(n2525), .A4(n2526), .ZN(n2522)
         );
  OAI221_X1 U2610 ( .B1(n169), .B2(n737), .C1(n393), .C2(n740), .A(n2527), 
        .ZN(n2526) );
  AOI22_X1 U2611 ( .A1(n743), .A2(n923), .B1(n746), .B2(n889), .ZN(n2527) );
  OAI221_X1 U2612 ( .B1(n170), .B2(n749), .C1(n394), .C2(n752), .A(n2528), 
        .ZN(n2525) );
  AOI22_X1 U2613 ( .A1(n755), .A2(n996), .B1(n758), .B2(n963), .ZN(n2528) );
  OAI221_X1 U2614 ( .B1(n171), .B2(n761), .C1(n395), .C2(n764), .A(n2529), 
        .ZN(n2524) );
  AOI22_X1 U2615 ( .A1(n767), .A2(n1065), .B1(n770), .B2(n1032), .ZN(n2529) );
  OAI221_X1 U2616 ( .B1(n172), .B2(n773), .C1(n396), .C2(n776), .A(n2530), 
        .ZN(n2523) );
  AOI22_X1 U2617 ( .A1(n779), .A2(n1134), .B1(n782), .B2(n1101), .ZN(n2530) );
  NOR4_X1 U2618 ( .A1(n2531), .A2(n2532), .A3(n2533), .A4(n2534), .ZN(n2521)
         );
  OAI221_X1 U2619 ( .B1(n4168), .B2(n785), .C1(n4169), .C2(n788), .A(n2535), 
        .ZN(n2534) );
  AOI22_X1 U2620 ( .A1(n791), .A2(n4170), .B1(n794), .B2(n4171), .ZN(n2535) );
  OAI221_X1 U2621 ( .B1(n173), .B2(n797), .C1(n397), .C2(n800), .A(n2536), 
        .ZN(n2533) );
  AOI22_X1 U2622 ( .A1(n803), .A2(n1310), .B1(n806), .B2(n1343), .ZN(n2536) );
  OAI221_X1 U2623 ( .B1(n174), .B2(n809), .C1(n398), .C2(n812), .A(n2537), 
        .ZN(n2532) );
  AOI22_X1 U2624 ( .A1(n815), .A2(n1171), .B1(n818), .B2(n1204), .ZN(n2537) );
  OAI221_X1 U2625 ( .B1(n175), .B2(n821), .C1(n399), .C2(n824), .A(n2538), 
        .ZN(n2531) );
  AOI22_X1 U2626 ( .A1(n827), .A2(n1241), .B1(n830), .B2(n1274), .ZN(n2538) );
  NAND2_X1 U2627 ( .A1(n2539), .A2(n2540), .ZN(OUT1[15]) );
  NOR4_X1 U2628 ( .A1(n2541), .A2(n2542), .A3(n2543), .A4(n2544), .ZN(n2540)
         );
  OAI221_X1 U2629 ( .B1(n176), .B2(n737), .C1(n400), .C2(n740), .A(n2545), 
        .ZN(n2544) );
  AOI22_X1 U2630 ( .A1(n743), .A2(n924), .B1(n746), .B2(n890), .ZN(n2545) );
  OAI221_X1 U2631 ( .B1(n177), .B2(n749), .C1(n401), .C2(n752), .A(n2546), 
        .ZN(n2543) );
  AOI22_X1 U2632 ( .A1(n755), .A2(n997), .B1(n758), .B2(n964), .ZN(n2546) );
  OAI221_X1 U2633 ( .B1(n178), .B2(n761), .C1(n402), .C2(n764), .A(n2547), 
        .ZN(n2542) );
  AOI22_X1 U2634 ( .A1(n767), .A2(n1066), .B1(n770), .B2(n1033), .ZN(n2547) );
  OAI221_X1 U2635 ( .B1(n179), .B2(n773), .C1(n403), .C2(n776), .A(n2548), 
        .ZN(n2541) );
  AOI22_X1 U2636 ( .A1(n779), .A2(n1135), .B1(n782), .B2(n1102), .ZN(n2548) );
  NOR4_X1 U2637 ( .A1(n2549), .A2(n2550), .A3(n2551), .A4(n2552), .ZN(n2539)
         );
  OAI221_X1 U2638 ( .B1(n4186), .B2(n785), .C1(n4187), .C2(n788), .A(n2553), 
        .ZN(n2552) );
  AOI22_X1 U2639 ( .A1(n791), .A2(n4188), .B1(n794), .B2(n4189), .ZN(n2553) );
  OAI221_X1 U2640 ( .B1(n180), .B2(n797), .C1(n404), .C2(n800), .A(n2554), 
        .ZN(n2551) );
  AOI22_X1 U2641 ( .A1(n803), .A2(n1311), .B1(n806), .B2(n1344), .ZN(n2554) );
  OAI221_X1 U2642 ( .B1(n181), .B2(n809), .C1(n405), .C2(n812), .A(n2555), 
        .ZN(n2550) );
  AOI22_X1 U2643 ( .A1(n815), .A2(n1172), .B1(n818), .B2(n1205), .ZN(n2555) );
  OAI221_X1 U2644 ( .B1(n182), .B2(n821), .C1(n406), .C2(n824), .A(n2556), 
        .ZN(n2549) );
  AOI22_X1 U2645 ( .A1(n827), .A2(n1242), .B1(n830), .B2(n1275), .ZN(n2556) );
  NAND2_X1 U2646 ( .A1(n2557), .A2(n2558), .ZN(OUT1[14]) );
  NOR4_X1 U2647 ( .A1(n2559), .A2(n2560), .A3(n2561), .A4(n2562), .ZN(n2558)
         );
  OAI221_X1 U2648 ( .B1(n183), .B2(n737), .C1(n407), .C2(n740), .A(n2563), 
        .ZN(n2562) );
  AOI22_X1 U2649 ( .A1(n743), .A2(n925), .B1(n746), .B2(n891), .ZN(n2563) );
  OAI221_X1 U2650 ( .B1(n184), .B2(n749), .C1(n408), .C2(n752), .A(n2564), 
        .ZN(n2561) );
  AOI22_X1 U2651 ( .A1(n755), .A2(n998), .B1(n758), .B2(n965), .ZN(n2564) );
  OAI221_X1 U2652 ( .B1(n185), .B2(n761), .C1(n409), .C2(n764), .A(n2565), 
        .ZN(n2560) );
  AOI22_X1 U2653 ( .A1(n767), .A2(n1067), .B1(n770), .B2(n1034), .ZN(n2565) );
  OAI221_X1 U2654 ( .B1(n186), .B2(n773), .C1(n410), .C2(n776), .A(n2566), 
        .ZN(n2559) );
  AOI22_X1 U2655 ( .A1(n779), .A2(n1136), .B1(n782), .B2(n1103), .ZN(n2566) );
  NOR4_X1 U2656 ( .A1(n2567), .A2(n2568), .A3(n2569), .A4(n2570), .ZN(n2557)
         );
  OAI221_X1 U2657 ( .B1(n4204), .B2(n785), .C1(n4205), .C2(n788), .A(n2571), 
        .ZN(n2570) );
  AOI22_X1 U2658 ( .A1(n791), .A2(n4206), .B1(n794), .B2(n4207), .ZN(n2571) );
  OAI221_X1 U2659 ( .B1(n187), .B2(n797), .C1(n411), .C2(n800), .A(n2572), 
        .ZN(n2569) );
  AOI22_X1 U2660 ( .A1(n803), .A2(n1312), .B1(n806), .B2(n1345), .ZN(n2572) );
  OAI221_X1 U2661 ( .B1(n188), .B2(n809), .C1(n412), .C2(n812), .A(n2573), 
        .ZN(n2568) );
  AOI22_X1 U2662 ( .A1(n815), .A2(n1173), .B1(n818), .B2(n1206), .ZN(n2573) );
  OAI221_X1 U2663 ( .B1(n189), .B2(n821), .C1(n413), .C2(n824), .A(n2574), 
        .ZN(n2567) );
  AOI22_X1 U2664 ( .A1(n827), .A2(n1243), .B1(n830), .B2(n1276), .ZN(n2574) );
  NAND2_X1 U2665 ( .A1(n2575), .A2(n2576), .ZN(OUT1[13]) );
  NOR4_X1 U2666 ( .A1(n2577), .A2(n2578), .A3(n2579), .A4(n2580), .ZN(n2576)
         );
  OAI221_X1 U2667 ( .B1(n190), .B2(n737), .C1(n414), .C2(n740), .A(n2581), 
        .ZN(n2580) );
  AOI22_X1 U2668 ( .A1(n743), .A2(n926), .B1(n746), .B2(n892), .ZN(n2581) );
  OAI221_X1 U2669 ( .B1(n191), .B2(n749), .C1(n415), .C2(n752), .A(n2582), 
        .ZN(n2579) );
  AOI22_X1 U2670 ( .A1(n755), .A2(n999), .B1(n758), .B2(n966), .ZN(n2582) );
  OAI221_X1 U2671 ( .B1(n192), .B2(n761), .C1(n416), .C2(n764), .A(n2583), 
        .ZN(n2578) );
  AOI22_X1 U2672 ( .A1(n767), .A2(n1068), .B1(n770), .B2(n1035), .ZN(n2583) );
  OAI221_X1 U2673 ( .B1(n193), .B2(n773), .C1(n417), .C2(n776), .A(n2584), 
        .ZN(n2577) );
  AOI22_X1 U2674 ( .A1(n779), .A2(n1137), .B1(n782), .B2(n1104), .ZN(n2584) );
  NOR4_X1 U2675 ( .A1(n2585), .A2(n2586), .A3(n2587), .A4(n2588), .ZN(n2575)
         );
  OAI221_X1 U2676 ( .B1(n4222), .B2(n785), .C1(n4223), .C2(n788), .A(n2589), 
        .ZN(n2588) );
  AOI22_X1 U2677 ( .A1(n791), .A2(n4224), .B1(n794), .B2(n4225), .ZN(n2589) );
  OAI221_X1 U2678 ( .B1(n194), .B2(n797), .C1(n418), .C2(n800), .A(n2590), 
        .ZN(n2587) );
  AOI22_X1 U2679 ( .A1(n803), .A2(n1313), .B1(n806), .B2(n1346), .ZN(n2590) );
  OAI221_X1 U2680 ( .B1(n195), .B2(n809), .C1(n419), .C2(n812), .A(n2591), 
        .ZN(n2586) );
  AOI22_X1 U2681 ( .A1(n815), .A2(n1174), .B1(n818), .B2(n1207), .ZN(n2591) );
  OAI221_X1 U2682 ( .B1(n196), .B2(n821), .C1(n420), .C2(n824), .A(n2592), 
        .ZN(n2585) );
  AOI22_X1 U2683 ( .A1(n827), .A2(n1244), .B1(n830), .B2(n1277), .ZN(n2592) );
  NAND2_X1 U2684 ( .A1(n2593), .A2(n2594), .ZN(OUT1[12]) );
  NOR4_X1 U2685 ( .A1(n2595), .A2(n2596), .A3(n2597), .A4(n2598), .ZN(n2594)
         );
  OAI221_X1 U2686 ( .B1(n197), .B2(n737), .C1(n421), .C2(n740), .A(n2599), 
        .ZN(n2598) );
  AOI22_X1 U2687 ( .A1(n743), .A2(n927), .B1(n746), .B2(n893), .ZN(n2599) );
  OAI221_X1 U2688 ( .B1(n198), .B2(n749), .C1(n422), .C2(n752), .A(n2600), 
        .ZN(n2597) );
  AOI22_X1 U2689 ( .A1(n755), .A2(n1000), .B1(n758), .B2(n967), .ZN(n2600) );
  OAI221_X1 U2690 ( .B1(n199), .B2(n761), .C1(n423), .C2(n764), .A(n2601), 
        .ZN(n2596) );
  AOI22_X1 U2691 ( .A1(n767), .A2(n1069), .B1(n770), .B2(n1036), .ZN(n2601) );
  OAI221_X1 U2692 ( .B1(n200), .B2(n773), .C1(n424), .C2(n776), .A(n2602), 
        .ZN(n2595) );
  AOI22_X1 U2693 ( .A1(n779), .A2(n1138), .B1(n782), .B2(n1105), .ZN(n2602) );
  NOR4_X1 U2694 ( .A1(n2603), .A2(n2604), .A3(n2605), .A4(n2606), .ZN(n2593)
         );
  OAI221_X1 U2695 ( .B1(n4240), .B2(n785), .C1(n4241), .C2(n788), .A(n2607), 
        .ZN(n2606) );
  AOI22_X1 U2696 ( .A1(n791), .A2(n4242), .B1(n794), .B2(n4243), .ZN(n2607) );
  OAI221_X1 U2697 ( .B1(n201), .B2(n797), .C1(n425), .C2(n800), .A(n2608), 
        .ZN(n2605) );
  AOI22_X1 U2698 ( .A1(n803), .A2(n1314), .B1(n806), .B2(n1347), .ZN(n2608) );
  OAI221_X1 U2699 ( .B1(n202), .B2(n809), .C1(n426), .C2(n812), .A(n2609), 
        .ZN(n2604) );
  AOI22_X1 U2700 ( .A1(n815), .A2(n1175), .B1(n818), .B2(n1208), .ZN(n2609) );
  OAI221_X1 U2701 ( .B1(n203), .B2(n821), .C1(n427), .C2(n824), .A(n2610), 
        .ZN(n2603) );
  AOI22_X1 U2702 ( .A1(n827), .A2(n1245), .B1(n830), .B2(n1278), .ZN(n2610) );
  NAND2_X1 U2703 ( .A1(n2611), .A2(n2612), .ZN(OUT1[11]) );
  NOR4_X1 U2704 ( .A1(n2613), .A2(n2614), .A3(n2615), .A4(n2616), .ZN(n2612)
         );
  OAI221_X1 U2705 ( .B1(n204), .B2(n737), .C1(n428), .C2(n740), .A(n2617), 
        .ZN(n2616) );
  AOI22_X1 U2706 ( .A1(n743), .A2(n928), .B1(n746), .B2(n894), .ZN(n2617) );
  OAI221_X1 U2707 ( .B1(n205), .B2(n749), .C1(n429), .C2(n752), .A(n2618), 
        .ZN(n2615) );
  AOI22_X1 U2708 ( .A1(n755), .A2(n1001), .B1(n758), .B2(n968), .ZN(n2618) );
  OAI221_X1 U2709 ( .B1(n206), .B2(n761), .C1(n430), .C2(n764), .A(n2619), 
        .ZN(n2614) );
  AOI22_X1 U2710 ( .A1(n767), .A2(n1070), .B1(n770), .B2(n1037), .ZN(n2619) );
  OAI221_X1 U2711 ( .B1(n207), .B2(n773), .C1(n431), .C2(n776), .A(n2620), 
        .ZN(n2613) );
  AOI22_X1 U2712 ( .A1(n779), .A2(n1139), .B1(n782), .B2(n1106), .ZN(n2620) );
  NOR4_X1 U2713 ( .A1(n2621), .A2(n2622), .A3(n2623), .A4(n2624), .ZN(n2611)
         );
  OAI221_X1 U2714 ( .B1(n4258), .B2(n785), .C1(n4259), .C2(n788), .A(n2625), 
        .ZN(n2624) );
  AOI22_X1 U2715 ( .A1(n791), .A2(n4260), .B1(n794), .B2(n4261), .ZN(n2625) );
  OAI221_X1 U2716 ( .B1(n208), .B2(n797), .C1(n432), .C2(n800), .A(n2626), 
        .ZN(n2623) );
  AOI22_X1 U2717 ( .A1(n803), .A2(n1315), .B1(n806), .B2(n1348), .ZN(n2626) );
  OAI221_X1 U2718 ( .B1(n209), .B2(n809), .C1(n433), .C2(n812), .A(n2627), 
        .ZN(n2622) );
  AOI22_X1 U2719 ( .A1(n815), .A2(n1176), .B1(n818), .B2(n1209), .ZN(n2627) );
  OAI221_X1 U2720 ( .B1(n210), .B2(n821), .C1(n434), .C2(n824), .A(n2628), 
        .ZN(n2621) );
  AOI22_X1 U2721 ( .A1(n827), .A2(n1246), .B1(n830), .B2(n1279), .ZN(n2628) );
  NAND2_X1 U2722 ( .A1(n2629), .A2(n2630), .ZN(OUT1[10]) );
  NOR4_X1 U2723 ( .A1(n2631), .A2(n2632), .A3(n2633), .A4(n2634), .ZN(n2630)
         );
  OAI221_X1 U2724 ( .B1(n211), .B2(n737), .C1(n435), .C2(n740), .A(n2635), 
        .ZN(n2634) );
  AOI22_X1 U2725 ( .A1(n743), .A2(n929), .B1(n746), .B2(n895), .ZN(n2635) );
  OAI221_X1 U2726 ( .B1(n212), .B2(n749), .C1(n436), .C2(n752), .A(n2636), 
        .ZN(n2633) );
  AOI22_X1 U2727 ( .A1(n755), .A2(n1002), .B1(n758), .B2(n969), .ZN(n2636) );
  OAI221_X1 U2728 ( .B1(n213), .B2(n761), .C1(n437), .C2(n764), .A(n2637), 
        .ZN(n2632) );
  AOI22_X1 U2729 ( .A1(n767), .A2(n1071), .B1(n770), .B2(n1038), .ZN(n2637) );
  OAI221_X1 U2730 ( .B1(n214), .B2(n773), .C1(n438), .C2(n776), .A(n2638), 
        .ZN(n2631) );
  AOI22_X1 U2731 ( .A1(n779), .A2(n1140), .B1(n782), .B2(n1107), .ZN(n2638) );
  NOR4_X1 U2732 ( .A1(n2639), .A2(n2640), .A3(n2641), .A4(n2642), .ZN(n2629)
         );
  OAI221_X1 U2733 ( .B1(n4276), .B2(n785), .C1(n4277), .C2(n788), .A(n2643), 
        .ZN(n2642) );
  AOI22_X1 U2734 ( .A1(n791), .A2(n4278), .B1(n794), .B2(n4279), .ZN(n2643) );
  OAI221_X1 U2735 ( .B1(n215), .B2(n797), .C1(n439), .C2(n800), .A(n2644), 
        .ZN(n2641) );
  AOI22_X1 U2736 ( .A1(n803), .A2(n1316), .B1(n806), .B2(n1349), .ZN(n2644) );
  OAI221_X1 U2737 ( .B1(n216), .B2(n809), .C1(n440), .C2(n812), .A(n2645), 
        .ZN(n2640) );
  AOI22_X1 U2738 ( .A1(n815), .A2(n1177), .B1(n818), .B2(n1210), .ZN(n2645) );
  OAI221_X1 U2739 ( .B1(n217), .B2(n821), .C1(n441), .C2(n824), .A(n2646), 
        .ZN(n2639) );
  AOI22_X1 U2740 ( .A1(n827), .A2(n1247), .B1(n830), .B2(n1280), .ZN(n2646) );
  NAND2_X1 U2741 ( .A1(n2647), .A2(n2648), .ZN(OUT1[0]) );
  NOR4_X1 U2742 ( .A1(n2649), .A2(n2650), .A3(n2651), .A4(n2652), .ZN(n2648)
         );
  OAI221_X1 U2743 ( .B1(n218), .B2(n737), .C1(n442), .C2(n740), .A(n2653), 
        .ZN(n2652) );
  AOI22_X1 U2744 ( .A1(n743), .A2(n939), .B1(n746), .B2(n905), .ZN(n2653) );
  AND2_X1 U2745 ( .A1(n2654), .A2(n2655), .ZN(n2067) );
  AND2_X1 U2746 ( .A1(n2656), .A2(n2655), .ZN(n2066) );
  NAND2_X1 U2747 ( .A1(n2654), .A2(n3682), .ZN(n2064) );
  NAND2_X1 U2748 ( .A1(n2656), .A2(n3682), .ZN(n2063) );
  OAI221_X1 U2749 ( .B1(n219), .B2(n749), .C1(n443), .C2(n752), .A(n3683), 
        .ZN(n2651) );
  AOI22_X1 U2750 ( .A1(n755), .A2(n1012), .B1(n758), .B2(n979), .ZN(n3683) );
  AND2_X1 U2751 ( .A1(n2654), .A2(n3684), .ZN(n2072) );
  AND2_X1 U2752 ( .A1(n2656), .A2(n3684), .ZN(n2071) );
  NAND2_X1 U2753 ( .A1(n2654), .A2(n3685), .ZN(n2069) );
  NOR3_X1 U2754 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n2654) );
  NAND2_X1 U2755 ( .A1(n2656), .A2(n3685), .ZN(n2068) );
  NOR3_X1 U2756 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n3686), .ZN(n2656) );
  OAI221_X1 U2757 ( .B1(n220), .B2(n761), .C1(n444), .C2(n764), .A(n3687), 
        .ZN(n2650) );
  AOI22_X1 U2758 ( .A1(n767), .A2(n1081), .B1(n770), .B2(n1048), .ZN(n3687) );
  AND2_X1 U2759 ( .A1(n2655), .A2(n3688), .ZN(n2077) );
  AND2_X1 U2760 ( .A1(n2655), .A2(n3689), .ZN(n2076) );
  NAND2_X1 U2761 ( .A1(n3682), .A2(n3688), .ZN(n2074) );
  NAND2_X1 U2762 ( .A1(n3682), .A2(n3689), .ZN(n2073) );
  OAI221_X1 U2763 ( .B1(n221), .B2(n773), .C1(n445), .C2(n776), .A(n3690), 
        .ZN(n2649) );
  AOI22_X1 U2764 ( .A1(n779), .A2(n1150), .B1(n782), .B2(n1117), .ZN(n3690) );
  AND2_X1 U2765 ( .A1(n3688), .A2(n3684), .ZN(n2082) );
  AND2_X1 U2766 ( .A1(n3689), .A2(n3684), .ZN(n2081) );
  NAND2_X1 U2767 ( .A1(n3685), .A2(n3688), .ZN(n2079) );
  NOR3_X1 U2768 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n3691), .ZN(n3688) );
  NAND2_X1 U2769 ( .A1(n3685), .A2(n3689), .ZN(n2078) );
  NOR3_X1 U2770 ( .A1(n3686), .A2(ADD_RD1[4]), .A3(n3691), .ZN(n3689) );
  NOR4_X1 U2771 ( .A1(n3692), .A2(n3693), .A3(n3694), .A4(n3695), .ZN(n2647)
         );
  OAI221_X1 U2772 ( .B1(n4294), .B2(n785), .C1(n4295), .C2(n788), .A(n3696), 
        .ZN(n3695) );
  AOI22_X1 U2773 ( .A1(n791), .A2(n4296), .B1(n794), .B2(n4297), .ZN(n3696) );
  AND2_X1 U2774 ( .A1(n3697), .A2(n3684), .ZN(n2091) );
  AND2_X1 U2775 ( .A1(n3698), .A2(n3684), .ZN(n2090) );
  NAND2_X1 U2776 ( .A1(n3698), .A2(n3685), .ZN(n2088) );
  NAND2_X1 U2777 ( .A1(n3697), .A2(n3685), .ZN(n2087) );
  OAI221_X1 U2778 ( .B1(n222), .B2(n797), .C1(n446), .C2(n800), .A(n3699), 
        .ZN(n3694) );
  AOI22_X1 U2779 ( .A1(n803), .A2(n1326), .B1(n806), .B2(n1359), .ZN(n3699) );
  AND2_X1 U2780 ( .A1(n3698), .A2(n2655), .ZN(n2096) );
  AND2_X1 U2781 ( .A1(n3697), .A2(n2655), .ZN(n2095) );
  NAND2_X1 U2782 ( .A1(n3697), .A2(n3682), .ZN(n2093) );
  NOR3_X1 U2783 ( .A1(n3691), .A2(ADD_RD1[0]), .A3(n3700), .ZN(n3697) );
  NAND2_X1 U2784 ( .A1(n3698), .A2(n3682), .ZN(n2092) );
  NOR3_X1 U2785 ( .A1(n3691), .A2(n3686), .A3(n3700), .ZN(n3698) );
  INV_X1 U2786 ( .A(ADD_RD1[3]), .ZN(n3691) );
  OAI221_X1 U2787 ( .B1(n223), .B2(n809), .C1(n447), .C2(n812), .A(n3701), 
        .ZN(n3693) );
  AOI22_X1 U2788 ( .A1(n815), .A2(n1187), .B1(n818), .B2(n1220), .ZN(n3701) );
  AND2_X1 U2789 ( .A1(n3702), .A2(n2655), .ZN(n2101) );
  AND2_X1 U2790 ( .A1(n3703), .A2(n2655), .ZN(n2100) );
  NOR3_X1 U2791 ( .A1(n3704), .A2(ADD_RD1[2]), .A3(n3705), .ZN(n2655) );
  NAND2_X1 U2792 ( .A1(n3702), .A2(n3682), .ZN(n2098) );
  NAND2_X1 U2793 ( .A1(n3703), .A2(n3682), .ZN(n2097) );
  OAI221_X1 U2794 ( .B1(n224), .B2(n821), .C1(n448), .C2(n824), .A(n3706), 
        .ZN(n3692) );
  AOI22_X1 U2795 ( .A1(n827), .A2(n1257), .B1(n830), .B2(n1290), .ZN(n3706) );
  AND2_X1 U2796 ( .A1(n3702), .A2(n3684), .ZN(n2106) );
  AND2_X1 U2797 ( .A1(n3703), .A2(n3684), .ZN(n2105) );
  NOR3_X1 U2798 ( .A1(n3707), .A2(n3704), .A3(n3705), .ZN(n3684) );
  NAND2_X1 U2799 ( .A1(n3702), .A2(n3685), .ZN(n2103) );
  NOR3_X1 U2800 ( .A1(n3686), .A2(ADD_RD1[3]), .A3(n3700), .ZN(n3702) );
  INV_X1 U2801 ( .A(ADD_RD1[0]), .ZN(n3686) );
  NAND2_X1 U2802 ( .A1(n3703), .A2(n3685), .ZN(n2102) );
  NOR3_X1 U2803 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n3700), .ZN(n3703) );
  AOI211_X1 U2804 ( .C1(n3708), .C2(n3709), .A(n1151), .B(n835), .ZN(N4192) );
  INV_X1 U2805 ( .A(WR), .ZN(n1151) );
  NAND4_X1 U2806 ( .A1(n3710), .A2(n3711), .A3(n3712), .A4(n3713), .ZN(n3709)
         );
  NOR3_X1 U2807 ( .A1(n3714), .A2(n3705), .A3(n3715), .ZN(n3713) );
  XOR2_X1 U2808 ( .A(ADD_WR[0]), .B(ADD_RD1[0]), .Z(n3715) );
  INV_X1 U2809 ( .A(RD1), .ZN(n3705) );
  XOR2_X1 U2810 ( .A(ADD_WR[3]), .B(ADD_RD1[3]), .Z(n3714) );
  XOR2_X1 U2811 ( .A(n3707), .B(ADD_WR[2]), .Z(n3712) );
  INV_X1 U2812 ( .A(ADD_RD1[2]), .ZN(n3707) );
  XOR2_X1 U2813 ( .A(ADD_WR[4]), .B(n3700), .Z(n3711) );
  INV_X1 U2814 ( .A(ADD_RD1[4]), .ZN(n3700) );
  XOR2_X1 U2815 ( .A(n3704), .B(ADD_WR[1]), .Z(n3710) );
  INV_X1 U2816 ( .A(ADD_RD1[1]), .ZN(n3704) );
  NAND4_X1 U2817 ( .A1(n3716), .A2(n3717), .A3(n3718), .A4(n3719), .ZN(n3708)
         );
  NOR3_X1 U2818 ( .A1(n3720), .A2(n2054), .A3(n3721), .ZN(n3719) );
  XOR2_X1 U2819 ( .A(ADD_WR[0]), .B(ADD_RD2[0]), .Z(n3721) );
  INV_X1 U2820 ( .A(RD2), .ZN(n2054) );
  XOR2_X1 U2821 ( .A(ADD_WR[3]), .B(ADD_RD2[3]), .Z(n3720) );
  XOR2_X1 U2822 ( .A(n2056), .B(ADD_WR[2]), .Z(n3718) );
  INV_X1 U2823 ( .A(ADD_RD2[2]), .ZN(n2056) );
  XOR2_X1 U2824 ( .A(ADD_WR[4]), .B(n2049), .Z(n3717) );
  INV_X1 U2825 ( .A(ADD_RD2[4]), .ZN(n2049) );
  XOR2_X1 U2826 ( .A(n2053), .B(ADD_WR[1]), .Z(n3716) );
  INV_X1 U2827 ( .A(ADD_RD2[1]), .ZN(n2053) );
endmodule


module FETCH_UNIT_NB32_LS5_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[31] , \carry[30] , \carry[29] , \carry[28] ,
         \carry[27] , \carry[26] , \carry[25] , \carry[24] , \carry[23] ,
         \carry[22] , \carry[21] , \carry[20] , \carry[19] , \carry[18] ,
         \carry[17] , \carry[16] , \carry[15] , \carry[14] , \carry[13] ,
         \carry[12] , \carry[11] , \carry[10] , \carry[9] , \carry[8] ,
         \carry[7] , \carry[6] , \carry[5] , \carry[4] , \carry[3] ;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  AND2_X1 U1 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  XOR2_X1 U2 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  XOR2_X1 U3 ( .A(A[31]), .B(\carry[31] ), .Z(SUM[31]) );
  AND2_X1 U4 ( .A1(\carry[30] ), .A2(A[30]), .ZN(\carry[31] ) );
  XOR2_X1 U5 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  AND2_X1 U6 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  XOR2_X1 U7 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  AND2_X1 U8 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  XOR2_X1 U9 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  AND2_X1 U10 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  XOR2_X1 U11 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  AND2_X1 U12 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  XOR2_X1 U13 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  AND2_X1 U14 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  XOR2_X1 U15 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  AND2_X1 U16 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  XOR2_X1 U17 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  AND2_X1 U18 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  XOR2_X1 U19 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  AND2_X1 U20 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  XOR2_X1 U21 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  AND2_X1 U22 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  XOR2_X1 U23 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  AND2_X1 U24 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  XOR2_X1 U25 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  AND2_X1 U26 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  XOR2_X1 U27 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  AND2_X1 U28 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  XOR2_X1 U29 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  AND2_X1 U30 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  XOR2_X1 U31 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  AND2_X1 U32 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  XOR2_X1 U33 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  AND2_X1 U34 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  XOR2_X1 U35 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  AND2_X1 U36 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  XOR2_X1 U37 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  AND2_X1 U38 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  XOR2_X1 U39 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  AND2_X1 U40 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  XOR2_X1 U41 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  AND2_X1 U42 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  XOR2_X1 U43 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  AND2_X1 U44 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  XOR2_X1 U45 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  AND2_X1 U46 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  XOR2_X1 U47 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  AND2_X1 U48 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  XOR2_X1 U49 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  AND2_X1 U50 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  XOR2_X1 U51 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  AND2_X1 U52 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  XOR2_X1 U53 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  AND2_X1 U54 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  XOR2_X1 U55 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  INV_X1 U56 ( .A(\carry[3] ), .ZN(SUM[2]) );
  AND2_X1 U57 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  XOR2_X1 U58 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
endmodule


module MUX21_generic_NB32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n44, n45, n46, n47, n48, n49, n50, n51;

  INV_X1 U1 ( .A(n10), .ZN(n1) );
  BUF_X1 U2 ( .A(n7), .Z(n9) );
  BUF_X1 U3 ( .A(n4), .Z(n8) );
  BUF_X1 U4 ( .A(n11), .Z(n7) );
  BUF_X1 U5 ( .A(n11), .Z(n2) );
  BUF_X1 U6 ( .A(n11), .Z(n10) );
  BUF_X1 U7 ( .A(n11), .Z(n3) );
  BUF_X1 U8 ( .A(n8), .Z(n6) );
  BUF_X1 U9 ( .A(n8), .Z(n5) );
  BUF_X1 U10 ( .A(n11), .Z(n4) );
  INV_X1 U11 ( .A(n49), .ZN(Y[7]) );
  AOI22_X1 U12 ( .A1(A[7]), .A2(SEL), .B1(B[7]), .B2(n2), .ZN(n49) );
  INV_X1 U13 ( .A(n25), .ZN(Y[21]) );
  INV_X1 U14 ( .A(n29), .ZN(Y[25]) );
  INV_X1 U15 ( .A(n33), .ZN(Y[29]) );
  INV_X1 U16 ( .A(n36), .ZN(Y[30]) );
  INV_X1 U17 ( .A(n13), .ZN(Y[10]) );
  AOI22_X1 U18 ( .A1(A[10]), .A2(SEL), .B1(B[10]), .B2(n9), .ZN(n13) );
  INV_X1 U19 ( .A(n14), .ZN(Y[11]) );
  AOI22_X1 U20 ( .A1(A[11]), .A2(SEL), .B1(B[11]), .B2(n9), .ZN(n14) );
  INV_X1 U21 ( .A(n15), .ZN(Y[12]) );
  AOI22_X1 U22 ( .A1(A[12]), .A2(SEL), .B1(B[12]), .B2(n9), .ZN(n15) );
  INV_X1 U23 ( .A(n16), .ZN(Y[13]) );
  AOI22_X1 U24 ( .A1(A[13]), .A2(SEL), .B1(B[13]), .B2(n8), .ZN(n16) );
  INV_X1 U25 ( .A(n17), .ZN(Y[14]) );
  AOI22_X1 U26 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(n8), .ZN(n17) );
  INV_X1 U27 ( .A(n47), .ZN(Y[5]) );
  AOI22_X1 U28 ( .A1(A[5]), .A2(n1), .B1(B[5]), .B2(n3), .ZN(n47) );
  INV_X1 U29 ( .A(n50), .ZN(Y[8]) );
  AOI22_X1 U30 ( .A1(A[8]), .A2(n1), .B1(B[8]), .B2(n2), .ZN(n50) );
  INV_X1 U31 ( .A(n19), .ZN(Y[16]) );
  AOI22_X1 U32 ( .A1(A[16]), .A2(SEL), .B1(B[16]), .B2(n8), .ZN(n19) );
  INV_X1 U33 ( .A(n20), .ZN(Y[17]) );
  AOI22_X1 U34 ( .A1(A[17]), .A2(SEL), .B1(B[17]), .B2(n7), .ZN(n20) );
  INV_X1 U35 ( .A(n21), .ZN(Y[18]) );
  AOI22_X1 U36 ( .A1(A[18]), .A2(SEL), .B1(B[18]), .B2(n7), .ZN(n21) );
  INV_X1 U37 ( .A(n22), .ZN(Y[19]) );
  AOI22_X1 U38 ( .A1(A[19]), .A2(SEL), .B1(B[19]), .B2(n7), .ZN(n22) );
  INV_X1 U39 ( .A(n24), .ZN(Y[20]) );
  AOI22_X1 U40 ( .A1(A[20]), .A2(n1), .B1(B[20]), .B2(n6), .ZN(n24) );
  INV_X1 U41 ( .A(n26), .ZN(Y[22]) );
  AOI22_X1 U42 ( .A1(A[22]), .A2(n1), .B1(B[22]), .B2(n6), .ZN(n26) );
  INV_X1 U43 ( .A(n27), .ZN(Y[23]) );
  AOI22_X1 U44 ( .A1(A[23]), .A2(n1), .B1(B[23]), .B2(n6), .ZN(n27) );
  INV_X1 U45 ( .A(n28), .ZN(Y[24]) );
  AOI22_X1 U46 ( .A1(A[24]), .A2(n1), .B1(B[24]), .B2(n5), .ZN(n28) );
  INV_X1 U47 ( .A(n30), .ZN(Y[26]) );
  AOI22_X1 U48 ( .A1(A[26]), .A2(n1), .B1(B[26]), .B2(n5), .ZN(n30) );
  INV_X1 U49 ( .A(n32), .ZN(Y[28]) );
  AOI22_X1 U50 ( .A1(A[28]), .A2(n1), .B1(B[28]), .B2(n4), .ZN(n32) );
  INV_X1 U51 ( .A(n31), .ZN(Y[27]) );
  INV_X1 U52 ( .A(n18), .ZN(Y[15]) );
  AOI22_X1 U53 ( .A1(A[15]), .A2(SEL), .B1(B[15]), .B2(n8), .ZN(n18) );
  INV_X1 U54 ( .A(n51), .ZN(Y[9]) );
  AOI22_X1 U55 ( .A1(SEL), .A2(A[9]), .B1(B[9]), .B2(n2), .ZN(n51) );
  INV_X1 U56 ( .A(n34), .ZN(Y[2]) );
  AOI22_X1 U57 ( .A1(A[2]), .A2(n1), .B1(B[2]), .B2(n4), .ZN(n34) );
  INV_X1 U58 ( .A(n46), .ZN(Y[4]) );
  AOI22_X1 U59 ( .A1(A[4]), .A2(n1), .B1(B[4]), .B2(n3), .ZN(n46) );
  INV_X1 U60 ( .A(n48), .ZN(Y[6]) );
  AOI22_X1 U61 ( .A1(A[6]), .A2(n1), .B1(B[6]), .B2(n2), .ZN(n48) );
  INV_X1 U62 ( .A(n45), .ZN(Y[3]) );
  AOI22_X1 U63 ( .A1(A[3]), .A2(n1), .B1(B[3]), .B2(n3), .ZN(n45) );
  INV_X1 U64 ( .A(SEL), .ZN(n11) );
  INV_X1 U65 ( .A(n12), .ZN(Y[0]) );
  AOI22_X1 U66 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n9), .ZN(n12) );
  INV_X1 U67 ( .A(n23), .ZN(Y[1]) );
  AOI22_X1 U68 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n23) );
  INV_X1 U69 ( .A(n44), .ZN(Y[31]) );
  AOI22_X1 U70 ( .A1(A[30]), .A2(n1), .B1(B[30]), .B2(n4), .ZN(n36) );
  AOI22_X1 U71 ( .A1(A[31]), .A2(n1), .B1(B[31]), .B2(n3), .ZN(n44) );
  AOI22_X1 U72 ( .A1(A[27]), .A2(n1), .B1(B[27]), .B2(n5), .ZN(n31) );
  AOI22_X1 U73 ( .A1(A[29]), .A2(n1), .B1(B[29]), .B2(n4), .ZN(n33) );
  AOI22_X1 U74 ( .A1(A[21]), .A2(n1), .B1(B[21]), .B2(n6), .ZN(n25) );
  AOI22_X1 U75 ( .A1(A[25]), .A2(n1), .B1(B[25]), .B2(n5), .ZN(n29) );
endmodule


module FD_NB32_4 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n33, n34, n35;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n35), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n35), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n34), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n34), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n34), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n34), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n33), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n33), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n33), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n33), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n33), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n33), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n33), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n33), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n33), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n33), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n33), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n33), .Q(Q[0]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n34), .Q(Q[15]) );
  BUF_X1 U3 ( .A(RESET), .Z(n33) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
endmodule


module MUX21_generic_NB32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5, n6, n8, n7;

  CLKBUF_X1 U3 ( .A(n8), .Z(n1) );
  CLKBUF_X1 U4 ( .A(n8), .Z(n2) );
  CLKBUF_X1 U5 ( .A(n6), .Z(n3) );
  CLKBUF_X1 U6 ( .A(n8), .Z(n4) );
  CLKBUF_X1 U8 ( .A(n8), .Z(n5) );
  MUX2_X1 U10 ( .A(B[1]), .B(A[1]), .S(n6), .Z(Y[1]) );
  MUX2_X1 U11 ( .A(B[0]), .B(A[0]), .S(n6), .Z(Y[0]) );
  MUX2_X1 U12 ( .A(B[2]), .B(A[2]), .S(n8), .Z(Y[2]) );
  MUX2_X1 U13 ( .A(B[3]), .B(A[3]), .S(n6), .Z(Y[3]) );
  MUX2_X1 U17 ( .A(B[7]), .B(A[7]), .S(n6), .Z(Y[7]) );
  MUX2_X1 U18 ( .A(B[8]), .B(A[8]), .S(n8), .Z(Y[8]) );
  MUX2_X1 U19 ( .A(B[9]), .B(A[9]), .S(n6), .Z(Y[9]) );
  MUX2_X1 U20 ( .A(B[10]), .B(A[10]), .S(n8), .Z(Y[10]) );
  MUX2_X1 U21 ( .A(B[11]), .B(A[11]), .S(n6), .Z(Y[11]) );
  MUX2_X1 U22 ( .A(B[12]), .B(A[12]), .S(n6), .Z(Y[12]) );
  MUX2_X1 U23 ( .A(B[13]), .B(A[13]), .S(n8), .Z(Y[13]) );
  MUX2_X1 U24 ( .A(B[14]), .B(A[14]), .S(n8), .Z(Y[14]) );
  MUX2_X1 U25 ( .A(B[16]), .B(A[16]), .S(n5), .Z(Y[16]) );
  MUX2_X1 U26 ( .A(B[17]), .B(A[17]), .S(n5), .Z(Y[17]) );
  MUX2_X1 U27 ( .A(B[18]), .B(A[18]), .S(n5), .Z(Y[18]) );
  MUX2_X1 U28 ( .A(B[19]), .B(A[19]), .S(n3), .Z(Y[19]) );
  MUX2_X1 U29 ( .A(B[20]), .B(A[20]), .S(n1), .Z(Y[20]) );
  MUX2_X1 U30 ( .A(B[21]), .B(A[21]), .S(n5), .Z(Y[21]) );
  MUX2_X1 U31 ( .A(B[22]), .B(A[22]), .S(n4), .Z(Y[22]) );
  MUX2_X1 U32 ( .A(B[23]), .B(A[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U33 ( .A(B[24]), .B(A[24]), .S(n5), .Z(Y[24]) );
  MUX2_X1 U34 ( .A(B[25]), .B(A[25]), .S(n5), .Z(Y[25]) );
  MUX2_X1 U35 ( .A(B[26]), .B(A[26]), .S(n5), .Z(Y[26]) );
  MUX2_X1 U36 ( .A(B[27]), .B(A[27]), .S(n6), .Z(Y[27]) );
  MUX2_X1 U37 ( .A(B[28]), .B(A[28]), .S(n5), .Z(Y[28]) );
  MUX2_X1 U38 ( .A(B[29]), .B(A[29]), .S(n6), .Z(Y[29]) );
  MUX2_X1 U39 ( .A(B[30]), .B(A[30]), .S(n6), .Z(Y[30]) );
  MUX2_X1 U40 ( .A(B[31]), .B(A[31]), .S(n8), .Z(Y[31]) );
  MUX2_X1 U14 ( .A(B[4]), .B(A[4]), .S(n8), .Z(Y[4]) );
  MUX2_X1 U16 ( .A(B[6]), .B(A[6]), .S(n7), .Z(Y[6]) );
  MUX2_X1 U15 ( .A(B[5]), .B(A[5]), .S(n7), .Z(Y[5]) );
  BUF_X2 U1 ( .A(SEL), .Z(n7) );
  MUX2_X1 U2 ( .A(B[15]), .B(A[15]), .S(n7), .Z(Y[15]) );
  CLKBUF_X3 U7 ( .A(SEL), .Z(n6) );
  CLKBUF_X3 U9 ( .A(SEL), .Z(n8) );
endmodule


module FD_NB32_5 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n33, n34, n35;

  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n34), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n34), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n34), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n33), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n33), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n33), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n33), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n33), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n33), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n33), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n33), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n33), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n33), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n33), .Q(Q[0]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n33), .Q(Q[1]) );
  DFFR_X2 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n35), .Q(Q[31]) );
  BUF_X1 U3 ( .A(RESET), .Z(n33) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
  DFFR_X2 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n34), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n35), .Q(Q[30]) );
endmodule


module BP_NB32_BP_LEN4_0 ( CLK, RST, EX_PC, CURR_PC, NEXT_PC, NEW_PC, INST, 
        MISS_HIT, PRED );
  input [31:0] EX_PC;
  input [31:0] CURR_PC;
  input [31:0] NEXT_PC;
  input [31:0] NEW_PC;
  input [31:0] INST;
  output [1:0] MISS_HIT;
  output [31:0] PRED;
  input CLK, RST;
  wire   INST_31, INST_30, INST_29, INST_28, INST_27, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, \PRED_TABLE[0][1] , \PRED_TABLE[0][0] ,
         \PRED_TABLE[1][1] , \PRED_TABLE[1][0] , \PRED_TABLE[2][1] ,
         \PRED_TABLE[2][0] , \PRED_TABLE[3][1] , \PRED_TABLE[3][0] ,
         \PRED_TABLE[4][1] , \PRED_TABLE[4][0] , \PRED_TABLE[5][1] ,
         \PRED_TABLE[5][0] , \PRED_TABLE[6][1] , \PRED_TABLE[6][0] ,
         \PRED_TABLE[7][1] , \PRED_TABLE[7][0] , \PRED_TABLE[8][1] ,
         \PRED_TABLE[8][0] , \PRED_TABLE[9][1] , \PRED_TABLE[9][0] ,
         \PRED_TABLE[10][1] , \PRED_TABLE[10][0] , \PRED_TABLE[11][1] ,
         \PRED_TABLE[11][0] , \PRED_TABLE[12][1] , \PRED_TABLE[12][0] ,
         \PRED_TABLE[13][1] , \PRED_TABLE[13][0] , \PRED_TABLE[14][1] ,
         \PRED_TABLE[14][0] , \PRED_TABLE[15][1] , \PRED_TABLE[15][0] ,
         \PRED_HISTORY[0][32] , \PRED_HISTORY[0][31] , \PRED_HISTORY[0][30] ,
         \PRED_HISTORY[0][29] , \PRED_HISTORY[0][28] , \PRED_HISTORY[0][27] ,
         \PRED_HISTORY[0][26] , \PRED_HISTORY[0][25] , \PRED_HISTORY[0][24] ,
         \PRED_HISTORY[0][23] , \PRED_HISTORY[0][22] , \PRED_HISTORY[0][21] ,
         \PRED_HISTORY[0][20] , \PRED_HISTORY[0][19] , \PRED_HISTORY[0][18] ,
         \PRED_HISTORY[0][17] , \PRED_HISTORY[0][16] , \PRED_HISTORY[0][15] ,
         \PRED_HISTORY[0][14] , \PRED_HISTORY[0][13] , \PRED_HISTORY[0][12] ,
         \PRED_HISTORY[0][11] , \PRED_HISTORY[0][10] , \PRED_HISTORY[0][9] ,
         \PRED_HISTORY[0][8] , \PRED_HISTORY[0][7] , \PRED_HISTORY[0][6] ,
         \PRED_HISTORY[0][5] , \PRED_HISTORY[0][4] , \PRED_HISTORY[0][3] ,
         \PRED_HISTORY[0][2] , \PRED_HISTORY[0][1] , \PRED_HISTORY[0][0] ,
         \PRED_HISTORY[1][31] , \PRED_HISTORY[1][30] , \PRED_HISTORY[1][29] ,
         \PRED_HISTORY[1][28] , \PRED_HISTORY[1][27] , \PRED_HISTORY[1][26] ,
         \PRED_HISTORY[1][25] , \PRED_HISTORY[1][24] , \PRED_HISTORY[1][23] ,
         \PRED_HISTORY[1][22] , \PRED_HISTORY[1][21] , \PRED_HISTORY[1][20] ,
         \PRED_HISTORY[1][19] , \PRED_HISTORY[1][18] , \PRED_HISTORY[1][17] ,
         \PRED_HISTORY[1][16] , \PRED_HISTORY[1][15] , \PRED_HISTORY[1][14] ,
         \PRED_HISTORY[1][13] , \PRED_HISTORY[1][12] , \PRED_HISTORY[1][11] ,
         \PRED_HISTORY[1][10] , \PRED_HISTORY[1][9] , \PRED_HISTORY[1][8] ,
         \PRED_HISTORY[1][7] , \PRED_HISTORY[1][6] , \PRED_HISTORY[1][5] ,
         \PRED_HISTORY[1][4] , \PRED_HISTORY[1][3] , \PRED_HISTORY[1][2] ,
         \PRED_HISTORY[1][1] , \PRED_HISTORY[1][0] , N815, \PC_HISTORY[0][3] ,
         \PC_HISTORY[0][2] , \PC_HISTORY[0][1] , \PC_HISTORY[0][0] ,
         \PC_HISTORY[1][3] , \PC_HISTORY[1][2] , \PC_HISTORY[1][1] ,
         \PC_HISTORY[1][0] , N849, N850, n8, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n45, n46, n47, n48,
         n49, n50, n51, n53, n54, n57, n60, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n90, n91, n93, n94, n95, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n135, n136, n174, n175, n176, n177, n180, n183, n186, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n387, n388, n390,
         n391, n393, n394, n396, n397, n398, n399, n400, n401, n404, n407,
         n408, n409, n413, n415, n417, n418, n419, n420, n424, n425, n426,
         n430, n431, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n863, n864, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n958, n959, n960, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n991, n992, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1055, n1056, n1057, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1119, n1120, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1150, n1151, n1152, n1153, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1183, n1184, n1185, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1214,
         n1215, n1216, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1247, n1248,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1360, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1476, n1477, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1571, n1572, n1573, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1604, n1605, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1668, n1669, n1670, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1732, n1733, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1763, n1764, n1765, n1766, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1796, n1797, n1798, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1827, n1828, n1829, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1860, n1861, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1, n2, n1963, n1964, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2218, n2219, n2220, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2366, n2321,
         n2320, n2319, n2237, n2221, n2217, n1965, n2367, n2368;
  wire   [31:0] PRED_TK;
  assign INST_31 = INST[31];
  assign INST_30 = INST[30];
  assign INST_29 = INST[29];
  assign INST_28 = INST[28];
  assign INST_27 = INST[27];

  DFFR_X1 \PRED_HISTORY_reg[0][32]  ( .D(n2330), .CK(CLK), .RN(n2205), .Q(
        \PRED_HISTORY[0][32] ) );
  DFFR_X1 \PC_HISTORY_reg[0][3]  ( .D(CURR_PC[5]), .CK(CLK), .RN(n2205), .Q(
        \PC_HISTORY[0][3] ) );
  DFFR_X1 \PC_HISTORY_reg[0][2]  ( .D(CURR_PC[4]), .CK(CLK), .RN(n2205), .Q(
        \PC_HISTORY[0][2] ) );
  DFFR_X1 \PC_HISTORY_reg[0][1]  ( .D(CURR_PC[3]), .CK(CLK), .RN(n2206), .Q(
        \PC_HISTORY[0][1] ) );
  DFFR_X1 \PC_HISTORY_reg[0][0]  ( .D(CURR_PC[2]), .CK(CLK), .RN(n2206), .Q(
        \PC_HISTORY[0][0] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][0]  ( .D(PRED[0]), .CK(CLK), .RN(n2206), .Q(
        \PRED_HISTORY[0][0] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][0]  ( .D(\PRED_HISTORY[0][0] ), .CK(CLK), .RN(
        n2206), .Q(\PRED_HISTORY[1][0] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][9]  ( .D(PRED[9]), .CK(CLK), .RN(n2206), .Q(
        \PRED_HISTORY[0][9] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][9]  ( .D(\PRED_HISTORY[0][9] ), .CK(CLK), .RN(
        n2206), .Q(\PRED_HISTORY[1][9] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][8]  ( .D(PRED[8]), .CK(CLK), .RN(n2206), .Q(
        \PRED_HISTORY[0][8] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][8]  ( .D(\PRED_HISTORY[0][8] ), .CK(CLK), .RN(
        n2207), .Q(\PRED_HISTORY[1][8] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][7]  ( .D(PRED[7]), .CK(CLK), .RN(n2207), .Q(
        \PRED_HISTORY[0][7] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][7]  ( .D(\PRED_HISTORY[0][7] ), .CK(CLK), .RN(
        n2207), .Q(\PRED_HISTORY[1][7] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][6]  ( .D(PRED[6]), .CK(CLK), .RN(n2207), .Q(
        \PRED_HISTORY[0][6] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][6]  ( .D(\PRED_HISTORY[0][6] ), .CK(CLK), .RN(
        n2207), .Q(\PRED_HISTORY[1][6] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][5]  ( .D(PRED[5]), .CK(CLK), .RN(n2207), .Q(
        \PRED_HISTORY[0][5] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][5]  ( .D(\PRED_HISTORY[0][5] ), .CK(CLK), .RN(
        n2207), .Q(\PRED_HISTORY[1][5] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][4]  ( .D(PRED[4]), .CK(CLK), .RN(n2207), .Q(
        \PRED_HISTORY[0][4] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][4]  ( .D(\PRED_HISTORY[0][4] ), .CK(CLK), .RN(
        n2207), .Q(\PRED_HISTORY[1][4] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][3]  ( .D(PRED[3]), .CK(CLK), .RN(n2207), .Q(
        \PRED_HISTORY[0][3] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][3]  ( .D(\PRED_HISTORY[0][3] ), .CK(CLK), .RN(
        n2207), .Q(\PRED_HISTORY[1][3] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][31]  ( .D(\PRED_HISTORY[0][31] ), .CK(CLK), 
        .RN(n2208), .Q(\PRED_HISTORY[1][31] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][30]  ( .D(\PRED_HISTORY[0][30] ), .CK(CLK), 
        .RN(n2208), .Q(\PRED_HISTORY[1][30] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][2]  ( .D(PRED[2]), .CK(CLK), .RN(n2208), .Q(
        \PRED_HISTORY[0][2] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][2]  ( .D(\PRED_HISTORY[0][2] ), .CK(CLK), .RN(
        n2208), .Q(\PRED_HISTORY[1][2] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][29]  ( .D(PRED[29]), .CK(CLK), .RN(n2208), .Q(
        \PRED_HISTORY[0][29] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][29]  ( .D(\PRED_HISTORY[0][29] ), .CK(CLK), 
        .RN(n2208), .Q(\PRED_HISTORY[1][29] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][28]  ( .D(PRED[28]), .CK(CLK), .RN(n2208), .Q(
        \PRED_HISTORY[0][28] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][28]  ( .D(\PRED_HISTORY[0][28] ), .CK(CLK), 
        .RN(n2208), .Q(\PRED_HISTORY[1][28] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][27]  ( .D(PRED[27]), .CK(CLK), .RN(n2208), .Q(
        \PRED_HISTORY[0][27] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][27]  ( .D(\PRED_HISTORY[0][27] ), .CK(CLK), 
        .RN(n2208), .Q(\PRED_HISTORY[1][27] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][26]  ( .D(PRED[26]), .CK(CLK), .RN(n2208), .Q(
        \PRED_HISTORY[0][26] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][26]  ( .D(\PRED_HISTORY[0][26] ), .CK(CLK), 
        .RN(n2209), .Q(\PRED_HISTORY[1][26] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][25]  ( .D(PRED[25]), .CK(CLK), .RN(n2209), .Q(
        \PRED_HISTORY[0][25] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][25]  ( .D(\PRED_HISTORY[0][25] ), .CK(CLK), 
        .RN(n2209), .Q(\PRED_HISTORY[1][25] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][24]  ( .D(PRED[24]), .CK(CLK), .RN(n2209), .Q(
        \PRED_HISTORY[0][24] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][24]  ( .D(\PRED_HISTORY[0][24] ), .CK(CLK), 
        .RN(n2209), .Q(\PRED_HISTORY[1][24] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][23]  ( .D(\PRED_HISTORY[0][23] ), .CK(CLK), 
        .RN(n2209), .Q(\PRED_HISTORY[1][23] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][22]  ( .D(PRED[22]), .CK(CLK), .RN(n2209), .Q(
        \PRED_HISTORY[0][22] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][22]  ( .D(\PRED_HISTORY[0][22] ), .CK(CLK), 
        .RN(n2209), .Q(\PRED_HISTORY[1][22] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][21]  ( .D(PRED[21]), .CK(CLK), .RN(n2209), .Q(
        \PRED_HISTORY[0][21] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][21]  ( .D(\PRED_HISTORY[0][21] ), .CK(CLK), 
        .RN(n2209), .Q(\PRED_HISTORY[1][21] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][20]  ( .D(PRED[20]), .CK(CLK), .RN(n2209), .Q(
        \PRED_HISTORY[0][20] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][20]  ( .D(\PRED_HISTORY[0][20] ), .CK(CLK), 
        .RN(n2210), .Q(\PRED_HISTORY[1][20] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][1]  ( .D(PRED[1]), .CK(CLK), .RN(n2210), .Q(
        \PRED_HISTORY[0][1] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][1]  ( .D(\PRED_HISTORY[0][1] ), .CK(CLK), .RN(
        n2210), .Q(\PRED_HISTORY[1][1] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][19]  ( .D(PRED[19]), .CK(CLK), .RN(n2210), .Q(
        \PRED_HISTORY[0][19] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][19]  ( .D(\PRED_HISTORY[0][19] ), .CK(CLK), 
        .RN(n2210), .Q(\PRED_HISTORY[1][19] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][18]  ( .D(PRED[18]), .CK(CLK), .RN(n2210), .Q(
        \PRED_HISTORY[0][18] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][18]  ( .D(\PRED_HISTORY[0][18] ), .CK(CLK), 
        .RN(n2210), .Q(\PRED_HISTORY[1][18] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][17]  ( .D(PRED[17]), .CK(CLK), .RN(n2210), .Q(
        \PRED_HISTORY[0][17] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][17]  ( .D(\PRED_HISTORY[0][17] ), .CK(CLK), 
        .RN(n2210), .Q(\PRED_HISTORY[1][17] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][16]  ( .D(PRED[16]), .CK(CLK), .RN(n2210), .Q(
        \PRED_HISTORY[0][16] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][16]  ( .D(\PRED_HISTORY[0][16] ), .CK(CLK), 
        .RN(n2210), .Q(\PRED_HISTORY[1][16] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][15]  ( .D(PRED[15]), .CK(CLK), .RN(n2210), .Q(
        \PRED_HISTORY[0][15] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][15]  ( .D(\PRED_HISTORY[0][15] ), .CK(CLK), 
        .RN(n2211), .Q(\PRED_HISTORY[1][15] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][14]  ( .D(PRED[14]), .CK(CLK), .RN(n2211), .Q(
        \PRED_HISTORY[0][14] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][14]  ( .D(\PRED_HISTORY[0][14] ), .CK(CLK), 
        .RN(n2211), .Q(\PRED_HISTORY[1][14] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][13]  ( .D(PRED[13]), .CK(CLK), .RN(n2211), .Q(
        \PRED_HISTORY[0][13] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][13]  ( .D(\PRED_HISTORY[0][13] ), .CK(CLK), 
        .RN(n2211), .Q(\PRED_HISTORY[1][13] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][12]  ( .D(PRED[12]), .CK(CLK), .RN(n2211), .Q(
        \PRED_HISTORY[0][12] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][12]  ( .D(\PRED_HISTORY[0][12] ), .CK(CLK), 
        .RN(n2211), .Q(\PRED_HISTORY[1][12] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][11]  ( .D(PRED[11]), .CK(CLK), .RN(n2211), .Q(
        \PRED_HISTORY[0][11] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][11]  ( .D(\PRED_HISTORY[0][11] ), .CK(CLK), 
        .RN(n2211), .Q(\PRED_HISTORY[1][11] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][10]  ( .D(PRED[10]), .CK(CLK), .RN(n2211), .Q(
        \PRED_HISTORY[0][10] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][10]  ( .D(\PRED_HISTORY[0][10] ), .CK(CLK), 
        .RN(n2211), .Q(\PRED_HISTORY[1][10] ) );
  DFFS_X1 \PRED_TABLE_reg[0][0]  ( .D(n1280), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[0][0] ), .QN(n731) );
  DFFS_X1 \PRED_TABLE_reg[2][0]  ( .D(n1279), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[2][0] ), .QN(n730) );
  DFFS_X1 \PRED_TABLE_reg[4][0]  ( .D(n1278), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[4][0] ), .QN(n729) );
  DFFS_X1 \PRED_TABLE_reg[6][0]  ( .D(n1277), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[6][0] ), .QN(n728) );
  DFFS_X1 \PRED_TABLE_reg[8][0]  ( .D(n1276), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[8][0] ), .QN(n727) );
  DFFS_X1 \PRED_TABLE_reg[10][0]  ( .D(n1275), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[10][0] ), .QN(n726) );
  DFFS_X1 \PRED_TABLE_reg[12][0]  ( .D(n1274), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[12][0] ), .QN(n725) );
  DFFS_X1 \PRED_TABLE_reg[14][0]  ( .D(n1273), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[14][0] ), .QN(n724) );
  DFFS_X1 \PRED_TABLE_reg[13][0]  ( .D(n1272), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[13][0] ), .QN(n723) );
  DFFS_X1 \PRED_TABLE_reg[11][0]  ( .D(n1271), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[11][0] ), .QN(n722) );
  DFFS_X1 \PRED_TABLE_reg[9][0]  ( .D(n1270), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[9][0] ), .QN(n721) );
  DFFS_X1 \PRED_TABLE_reg[7][0]  ( .D(n1269), .CK(CLK), .SN(n2212), .Q(
        \PRED_TABLE[7][0] ), .QN(n720) );
  DFFS_X1 \PRED_TABLE_reg[5][0]  ( .D(n1268), .CK(CLK), .SN(n2213), .Q(
        \PRED_TABLE[5][0] ), .QN(n719) );
  DFFS_X1 \PRED_TABLE_reg[3][0]  ( .D(n1267), .CK(CLK), .SN(n2213), .Q(
        \PRED_TABLE[3][0] ), .QN(n718) );
  DFFS_X1 \PRED_TABLE_reg[1][0]  ( .D(n1266), .CK(CLK), .SN(n2213), .Q(
        \PRED_TABLE[1][0] ), .QN(n717) );
  DFFS_X1 \PRED_TABLE_reg[15][0]  ( .D(n1265), .CK(CLK), .SN(n2213), .Q(
        \PRED_TABLE[15][0] ), .QN(n716) );
  DFFR_X1 \PC_TABLE_reg[9][5]  ( .D(n1575), .CK(CLK), .RN(RST), .Q(n444), .QN(
        n962) );
  DFFR_X1 \PC_TABLE_reg[8][5]  ( .D(n1607), .CK(CLK), .RN(RST), .Q(n443), .QN(
        n994) );
  DFFR_X1 \PC_TABLE_reg[5][2]  ( .D(n1699), .CK(CLK), .RN(RST), .Q(n387), .QN(
        n1086) );
  DFFR_X1 \PC_TABLE_reg[4][4]  ( .D(n1730), .CK(CLK), .RN(RST), .Q(n418), .QN(
        n1117) );
  DFFR_X1 \PC_TABLE_reg[1][2]  ( .D(n1827), .CK(CLK), .RN(RST), .Q(n390), .QN(
        n1214) );
  DFFR_X1 \PC_TABLE_reg[9][2]  ( .D(n1571), .CK(CLK), .RN(RST), .Q(n396), .QN(
        n958) );
  DFFR_X1 \PC_TABLE_reg[5][4]  ( .D(n1698), .CK(CLK), .RN(RST), .Q(n419), .QN(
        n1085) );
  DFFR_X1 \PC_TABLE_reg[2][3]  ( .D(n1798), .CK(CLK), .RN(RST), .QN(n1185) );
  DFFR_X1 \PC_TABLE_reg[6][4]  ( .D(n1666), .CK(CLK), .RN(RST), .QN(n1053) );
  DFFR_X1 \PC_TABLE_reg[6][3]  ( .D(n1670), .CK(CLK), .RN(RST), .QN(n1057) );
  DFFR_X1 \PC_TABLE_reg[12][5]  ( .D(n1479), .CK(CLK), .RN(RST), .QN(n866) );
  DFFR_X1 \PC_TABLE_reg[12][4]  ( .D(n1474), .CK(CLK), .RN(RST), .QN(n861) );
  DFFR_X1 \PC_TABLE_reg[7][4]  ( .D(n1634), .CK(CLK), .RN(RST), .QN(n1021) );
  DFFR_X1 \PC_TABLE_reg[7][3]  ( .D(n1638), .CK(CLK), .RN(RST), .QN(n1025) );
  DFFR_X1 \PC_TABLE_reg[7][2]  ( .D(n1635), .CK(CLK), .RN(RST), .QN(n1022) );
  DFFR_X1 \PC_TABLE_reg[10][5]  ( .D(n1543), .CK(CLK), .RN(RST), .QN(n930) );
  DFFR_X1 \PC_TABLE_reg[10][3]  ( .D(n1542), .CK(CLK), .RN(RST), .QN(n929) );
  DFFR_X1 \PC_TABLE_reg[3][3]  ( .D(n1766), .CK(CLK), .RN(RST), .QN(n1153) );
  DFFR_X1 \PC_TABLE_reg[3][2]  ( .D(n1763), .CK(CLK), .RN(RST), .QN(n1150) );
  DFFR_X1 \PC_TABLE_reg[13][5]  ( .D(n1447), .CK(CLK), .RN(RST), .QN(n834) );
  DFFR_X1 \PC_TABLE_reg[13][4]  ( .D(n1442), .CK(CLK), .RN(RST), .QN(n829) );
  DFFR_X1 \PC_TABLE_reg[13][2]  ( .D(n1443), .CK(CLK), .RN(RST), .QN(n830) );
  DFFR_X1 \PC_TABLE_reg[11][5]  ( .D(n1511), .CK(CLK), .RN(RST), .QN(n898) );
  DFFR_X1 \PC_TABLE_reg[11][3]  ( .D(n1510), .CK(CLK), .RN(RST), .QN(n897) );
  DFFR_X1 \PC_TABLE_reg[11][2]  ( .D(n1507), .CK(CLK), .RN(RST), .QN(n894) );
  DFFR_X1 \PC_TABLE_reg[2][27]  ( .D(n1810), .CK(CLK), .RN(RST), .QN(n1197) );
  DFFR_X1 \PC_TABLE_reg[2][25]  ( .D(n1809), .CK(CLK), .RN(RST), .QN(n1196) );
  DFFR_X1 \PC_TABLE_reg[2][23]  ( .D(n1808), .CK(CLK), .RN(RST), .QN(n1195) );
  DFFR_X1 \PC_TABLE_reg[2][21]  ( .D(n1807), .CK(CLK), .RN(RST), .QN(n1194) );
  DFFR_X1 \PC_TABLE_reg[6][26]  ( .D(n1655), .CK(CLK), .RN(RST), .QN(n1042) );
  DFFR_X1 \PC_TABLE_reg[6][24]  ( .D(n1656), .CK(CLK), .RN(RST), .QN(n1043) );
  DFFR_X1 \PC_TABLE_reg[6][22]  ( .D(n1657), .CK(CLK), .RN(RST), .QN(n1044) );
  DFFR_X1 \PC_TABLE_reg[6][20]  ( .D(n1658), .CK(CLK), .RN(RST), .QN(n1045) );
  DFFR_X1 \PC_TABLE_reg[12][26]  ( .D(n1463), .CK(CLK), .RN(RST), .QN(n850) );
  DFFR_X1 \PC_TABLE_reg[12][24]  ( .D(n1464), .CK(CLK), .RN(RST), .QN(n851) );
  DFFR_X1 \PC_TABLE_reg[12][22]  ( .D(n1465), .CK(CLK), .RN(RST), .QN(n852) );
  DFFR_X1 \PC_TABLE_reg[12][20]  ( .D(n1466), .CK(CLK), .RN(RST), .QN(n853) );
  DFFR_X1 \PC_TABLE_reg[2][28]  ( .D(n1782), .CK(CLK), .RN(RST), .QN(n1169) );
  DFFR_X1 \PC_TABLE_reg[2][26]  ( .D(n1783), .CK(CLK), .RN(RST), .QN(n1170) );
  DFFR_X1 \PC_TABLE_reg[2][24]  ( .D(n1784), .CK(CLK), .RN(RST), .QN(n1171) );
  DFFR_X1 \PC_TABLE_reg[2][19]  ( .D(n1806), .CK(CLK), .RN(RST), .QN(n1193) );
  DFFR_X1 \PC_TABLE_reg[2][17]  ( .D(n1805), .CK(CLK), .RN(RST), .QN(n1192) );
  DFFR_X1 \PC_TABLE_reg[2][15]  ( .D(n1804), .CK(CLK), .RN(RST), .QN(n1191) );
  DFFR_X1 \PC_TABLE_reg[2][10]  ( .D(n1791), .CK(CLK), .RN(RST), .QN(n1178) );
  DFFR_X1 \PC_TABLE_reg[2][8]  ( .D(n1792), .CK(CLK), .RN(RST), .QN(n1179) );
  DFFR_X1 \PC_TABLE_reg[2][6]  ( .D(n1793), .CK(CLK), .RN(RST), .QN(n1180) );
  DFFR_X1 \PC_TABLE_reg[2][31]  ( .D(n1812), .CK(CLK), .RN(RST), .QN(n1199) );
  DFFR_X1 \PC_TABLE_reg[2][30]  ( .D(n1781), .CK(CLK), .RN(RST), .QN(n1168) );
  DFFR_X1 \PC_TABLE_reg[2][29]  ( .D(n1811), .CK(CLK), .RN(RST), .QN(n1198) );
  DFFR_X1 \PC_TABLE_reg[2][16]  ( .D(n1788), .CK(CLK), .RN(RST), .QN(n1175) );
  DFFR_X1 \PC_TABLE_reg[2][14]  ( .D(n1789), .CK(CLK), .RN(RST), .QN(n1176) );
  DFFR_X1 \PC_TABLE_reg[2][13]  ( .D(n1803), .CK(CLK), .RN(RST), .QN(n1190) );
  DFFR_X1 \PC_TABLE_reg[2][12]  ( .D(n1790), .CK(CLK), .RN(RST), .QN(n1177) );
  DFFR_X1 \PC_TABLE_reg[2][11]  ( .D(n1802), .CK(CLK), .RN(RST), .QN(n1189) );
  DFFR_X1 \PC_TABLE_reg[2][9]  ( .D(n1801), .CK(CLK), .RN(RST), .QN(n1188) );
  DFFR_X1 \PC_TABLE_reg[7][25]  ( .D(n1649), .CK(CLK), .RN(RST), .QN(n1036) );
  DFFR_X1 \PC_TABLE_reg[7][21]  ( .D(n1647), .CK(CLK), .RN(RST), .QN(n1034) );
  DFFR_X1 \PC_TABLE_reg[7][14]  ( .D(n1629), .CK(CLK), .RN(RST), .QN(n1016) );
  DFFR_X1 \PC_TABLE_reg[7][7]  ( .D(n1640), .CK(CLK), .RN(RST), .QN(n1027) );
  DFFR_X1 \PC_TABLE_reg[7][1]  ( .D(n1637), .CK(CLK), .RN(RST), .QN(n1024) );
  DFFR_X1 \PC_TABLE_reg[7][30]  ( .D(n1621), .CK(CLK), .RN(RST), .QN(n1008) );
  DFFR_X1 \PC_TABLE_reg[7][29]  ( .D(n1651), .CK(CLK), .RN(RST), .QN(n1038) );
  DFFR_X1 \PC_TABLE_reg[7][23]  ( .D(n1648), .CK(CLK), .RN(RST), .QN(n1035) );
  DFFR_X1 \PC_TABLE_reg[7][16]  ( .D(n1628), .CK(CLK), .RN(RST), .QN(n1015) );
  DFFR_X1 \PC_TABLE_reg[7][13]  ( .D(n1643), .CK(CLK), .RN(RST), .QN(n1030) );
  DFFR_X1 \PC_TABLE_reg[7][10]  ( .D(n1631), .CK(CLK), .RN(RST), .QN(n1018) );
  DFFR_X1 \PC_TABLE_reg[7][9]  ( .D(n1641), .CK(CLK), .RN(RST), .QN(n1028) );
  DFFR_X1 \PC_TABLE_reg[7][31]  ( .D(n1652), .CK(CLK), .RN(RST), .QN(n1039) );
  DFFR_X1 \PC_TABLE_reg[7][28]  ( .D(n1622), .CK(CLK), .RN(RST), .QN(n1009) );
  DFFR_X1 \PC_TABLE_reg[7][27]  ( .D(n1650), .CK(CLK), .RN(RST), .QN(n1037) );
  DFFR_X1 \PC_TABLE_reg[7][20]  ( .D(n1626), .CK(CLK), .RN(RST), .QN(n1013) );
  DFFR_X1 \PC_TABLE_reg[7][19]  ( .D(n1646), .CK(CLK), .RN(RST), .QN(n1033) );
  DFFR_X1 \PC_TABLE_reg[7][17]  ( .D(n1645), .CK(CLK), .RN(RST), .QN(n1032) );
  DFFR_X1 \PC_TABLE_reg[7][15]  ( .D(n1644), .CK(CLK), .RN(RST), .QN(n1031) );
  DFFR_X1 \PC_TABLE_reg[7][12]  ( .D(n1630), .CK(CLK), .RN(RST), .QN(n1017) );
  DFFR_X1 \PC_TABLE_reg[7][11]  ( .D(n1642), .CK(CLK), .RN(RST), .QN(n1029) );
  DFFR_X1 \PC_TABLE_reg[7][8]  ( .D(n1632), .CK(CLK), .RN(RST), .QN(n1019) );
  DFFR_X1 \PC_TABLE_reg[7][6]  ( .D(n1633), .CK(CLK), .RN(RST), .QN(n1020) );
  DFFR_X1 \PC_TABLE_reg[7][0]  ( .D(n1636), .CK(CLK), .RN(RST), .QN(n1023) );
  DFFR_X1 \PC_TABLE_reg[2][22]  ( .D(n1785), .CK(CLK), .RN(RST), .QN(n1172) );
  DFFR_X1 \PC_TABLE_reg[2][20]  ( .D(n1786), .CK(CLK), .RN(RST), .QN(n1173) );
  DFFR_X1 \PC_TABLE_reg[2][18]  ( .D(n1787), .CK(CLK), .RN(RST), .QN(n1174) );
  DFFR_X1 \PC_TABLE_reg[2][7]  ( .D(n1800), .CK(CLK), .RN(RST), .QN(n1187) );
  DFFR_X1 \PC_TABLE_reg[2][1]  ( .D(n1797), .CK(CLK), .RN(RST), .QN(n1184) );
  DFFR_X1 \PC_TABLE_reg[2][0]  ( .D(n1796), .CK(CLK), .RN(RST), .QN(n1183) );
  DFFR_X1 \PC_TABLE_reg[6][28]  ( .D(n1654), .CK(CLK), .RN(RST), .QN(n1041) );
  DFFR_X1 \PC_TABLE_reg[6][27]  ( .D(n1682), .CK(CLK), .RN(RST), .QN(n1069) );
  DFFR_X1 \PC_TABLE_reg[6][12]  ( .D(n1662), .CK(CLK), .RN(RST), .QN(n1049) );
  DFFR_X1 \PC_TABLE_reg[6][11]  ( .D(n1674), .CK(CLK), .RN(RST), .QN(n1061) );
  DFFR_X1 \PC_TABLE_reg[6][7]  ( .D(n1672), .CK(CLK), .RN(RST), .QN(n1059) );
  DFFR_X1 \PC_TABLE_reg[6][1]  ( .D(n1669), .CK(CLK), .RN(RST), .QN(n1056) );
  DFFR_X1 \PC_TABLE_reg[6][31]  ( .D(n1684), .CK(CLK), .RN(RST), .QN(n1071) );
  DFFR_X1 \PC_TABLE_reg[6][30]  ( .D(n1653), .CK(CLK), .RN(RST), .QN(n1040) );
  DFFR_X1 \PC_TABLE_reg[6][29]  ( .D(n1683), .CK(CLK), .RN(RST), .QN(n1070) );
  DFFR_X1 \PC_TABLE_reg[6][25]  ( .D(n1681), .CK(CLK), .RN(RST), .QN(n1068) );
  DFFR_X1 \PC_TABLE_reg[6][14]  ( .D(n1661), .CK(CLK), .RN(RST), .QN(n1048) );
  DFFR_X1 \PC_TABLE_reg[6][10]  ( .D(n1663), .CK(CLK), .RN(RST), .QN(n1050) );
  DFFR_X1 \PC_TABLE_reg[6][9]  ( .D(n1673), .CK(CLK), .RN(RST), .QN(n1060) );
  DFFR_X1 \PC_TABLE_reg[6][8]  ( .D(n1664), .CK(CLK), .RN(RST), .QN(n1051) );
  DFFR_X1 \PC_TABLE_reg[13][25]  ( .D(n1457), .CK(CLK), .RN(RST), .QN(n844) );
  DFFR_X1 \PC_TABLE_reg[13][21]  ( .D(n1455), .CK(CLK), .RN(RST), .QN(n842) );
  DFFR_X1 \PC_TABLE_reg[13][14]  ( .D(n1437), .CK(CLK), .RN(RST), .QN(n824) );
  DFFR_X1 \PC_TABLE_reg[13][7]  ( .D(n1448), .CK(CLK), .RN(RST), .QN(n835) );
  DFFR_X1 \PC_TABLE_reg[13][1]  ( .D(n1445), .CK(CLK), .RN(RST), .QN(n832) );
  DFFR_X1 \PC_TABLE_reg[12][28]  ( .D(n1462), .CK(CLK), .RN(RST), .QN(n849) );
  DFFR_X1 \PC_TABLE_reg[12][27]  ( .D(n1490), .CK(CLK), .RN(RST), .QN(n877) );
  DFFR_X1 \PC_TABLE_reg[12][12]  ( .D(n1470), .CK(CLK), .RN(RST), .QN(n857) );
  DFFR_X1 \PC_TABLE_reg[12][11]  ( .D(n1482), .CK(CLK), .RN(RST), .QN(n869) );
  DFFR_X1 \PC_TABLE_reg[12][7]  ( .D(n1480), .CK(CLK), .RN(RST), .QN(n867) );
  DFFR_X1 \PC_TABLE_reg[12][1]  ( .D(n1477), .CK(CLK), .RN(RST), .QN(n864) );
  DFFR_X1 \PC_TABLE_reg[11][25]  ( .D(n1521), .CK(CLK), .RN(RST), .QN(n908) );
  DFFR_X1 \PC_TABLE_reg[11][21]  ( .D(n1519), .CK(CLK), .RN(RST), .QN(n906) );
  DFFR_X1 \PC_TABLE_reg[11][14]  ( .D(n1501), .CK(CLK), .RN(RST), .QN(n888) );
  DFFR_X1 \PC_TABLE_reg[11][7]  ( .D(n1512), .CK(CLK), .RN(RST), .QN(n899) );
  DFFR_X1 \PC_TABLE_reg[11][1]  ( .D(n1509), .CK(CLK), .RN(RST), .QN(n896) );
  DFFR_X1 \PC_TABLE_reg[13][30]  ( .D(n1429), .CK(CLK), .RN(RST), .QN(n816) );
  DFFR_X1 \PC_TABLE_reg[13][29]  ( .D(n1459), .CK(CLK), .RN(RST), .QN(n846) );
  DFFR_X1 \PC_TABLE_reg[13][23]  ( .D(n1456), .CK(CLK), .RN(RST), .QN(n843) );
  DFFR_X1 \PC_TABLE_reg[13][16]  ( .D(n1436), .CK(CLK), .RN(RST), .QN(n823) );
  DFFR_X1 \PC_TABLE_reg[13][13]  ( .D(n1451), .CK(CLK), .RN(RST), .QN(n838) );
  DFFR_X1 \PC_TABLE_reg[13][10]  ( .D(n1439), .CK(CLK), .RN(RST), .QN(n826) );
  DFFR_X1 \PC_TABLE_reg[13][9]  ( .D(n1449), .CK(CLK), .RN(RST), .QN(n836) );
  DFFR_X1 \PC_TABLE_reg[12][31]  ( .D(n1492), .CK(CLK), .RN(RST), .QN(n879) );
  DFFR_X1 \PC_TABLE_reg[12][30]  ( .D(n1461), .CK(CLK), .RN(RST), .QN(n848) );
  DFFR_X1 \PC_TABLE_reg[12][29]  ( .D(n1491), .CK(CLK), .RN(RST), .QN(n878) );
  DFFR_X1 \PC_TABLE_reg[12][25]  ( .D(n1489), .CK(CLK), .RN(RST), .QN(n876) );
  DFFR_X1 \PC_TABLE_reg[12][14]  ( .D(n1469), .CK(CLK), .RN(RST), .QN(n856) );
  DFFR_X1 \PC_TABLE_reg[12][10]  ( .D(n1471), .CK(CLK), .RN(RST), .QN(n858) );
  DFFR_X1 \PC_TABLE_reg[12][9]  ( .D(n1481), .CK(CLK), .RN(RST), .QN(n868) );
  DFFR_X1 \PC_TABLE_reg[12][8]  ( .D(n1472), .CK(CLK), .RN(RST), .QN(n859) );
  DFFR_X1 \PC_TABLE_reg[11][30]  ( .D(n1493), .CK(CLK), .RN(RST), .QN(n880) );
  DFFR_X1 \PC_TABLE_reg[11][29]  ( .D(n1523), .CK(CLK), .RN(RST), .QN(n910) );
  DFFR_X1 \PC_TABLE_reg[11][23]  ( .D(n1520), .CK(CLK), .RN(RST), .QN(n907) );
  DFFR_X1 \PC_TABLE_reg[11][16]  ( .D(n1500), .CK(CLK), .RN(RST), .QN(n887) );
  DFFR_X1 \PC_TABLE_reg[11][13]  ( .D(n1515), .CK(CLK), .RN(RST), .QN(n902) );
  DFFR_X1 \PC_TABLE_reg[11][10]  ( .D(n1503), .CK(CLK), .RN(RST), .QN(n890) );
  DFFR_X1 \PC_TABLE_reg[11][9]  ( .D(n1513), .CK(CLK), .RN(RST), .QN(n900) );
  DFFR_X1 \PC_TABLE_reg[6][23]  ( .D(n1680), .CK(CLK), .RN(RST), .QN(n1067) );
  DFFR_X1 \PC_TABLE_reg[6][21]  ( .D(n1679), .CK(CLK), .RN(RST), .QN(n1066) );
  DFFR_X1 \PC_TABLE_reg[6][19]  ( .D(n1678), .CK(CLK), .RN(RST), .QN(n1065) );
  DFFR_X1 \PC_TABLE_reg[6][18]  ( .D(n1659), .CK(CLK), .RN(RST), .QN(n1046) );
  DFFR_X1 \PC_TABLE_reg[6][17]  ( .D(n1677), .CK(CLK), .RN(RST), .QN(n1064) );
  DFFR_X1 \PC_TABLE_reg[6][16]  ( .D(n1660), .CK(CLK), .RN(RST), .QN(n1047) );
  DFFR_X1 \PC_TABLE_reg[6][15]  ( .D(n1676), .CK(CLK), .RN(RST), .QN(n1063) );
  DFFR_X1 \PC_TABLE_reg[6][13]  ( .D(n1675), .CK(CLK), .RN(RST), .QN(n1062) );
  DFFR_X1 \PC_TABLE_reg[6][6]  ( .D(n1665), .CK(CLK), .RN(RST), .QN(n1052) );
  DFFR_X1 \PC_TABLE_reg[6][0]  ( .D(n1668), .CK(CLK), .RN(RST), .QN(n1055) );
  DFFR_X1 \PC_TABLE_reg[13][31]  ( .D(n1460), .CK(CLK), .RN(RST), .QN(n847) );
  DFFR_X1 \PC_TABLE_reg[13][28]  ( .D(n1430), .CK(CLK), .RN(RST), .QN(n817) );
  DFFR_X1 \PC_TABLE_reg[13][27]  ( .D(n1458), .CK(CLK), .RN(RST), .QN(n845) );
  DFFR_X1 \PC_TABLE_reg[13][20]  ( .D(n1434), .CK(CLK), .RN(RST), .QN(n821) );
  DFFR_X1 \PC_TABLE_reg[13][19]  ( .D(n1454), .CK(CLK), .RN(RST), .QN(n841) );
  DFFR_X1 \PC_TABLE_reg[13][17]  ( .D(n1453), .CK(CLK), .RN(RST), .QN(n840) );
  DFFR_X1 \PC_TABLE_reg[13][15]  ( .D(n1452), .CK(CLK), .RN(RST), .QN(n839) );
  DFFR_X1 \PC_TABLE_reg[13][12]  ( .D(n1438), .CK(CLK), .RN(RST), .QN(n825) );
  DFFR_X1 \PC_TABLE_reg[13][11]  ( .D(n1450), .CK(CLK), .RN(RST), .QN(n837) );
  DFFR_X1 \PC_TABLE_reg[13][8]  ( .D(n1440), .CK(CLK), .RN(RST), .QN(n827) );
  DFFR_X1 \PC_TABLE_reg[13][6]  ( .D(n1441), .CK(CLK), .RN(RST), .QN(n828) );
  DFFR_X1 \PC_TABLE_reg[13][0]  ( .D(n1444), .CK(CLK), .RN(RST), .QN(n831) );
  DFFR_X1 \PC_TABLE_reg[12][23]  ( .D(n1488), .CK(CLK), .RN(RST), .QN(n875) );
  DFFR_X1 \PC_TABLE_reg[12][21]  ( .D(n1487), .CK(CLK), .RN(RST), .QN(n874) );
  DFFR_X1 \PC_TABLE_reg[12][19]  ( .D(n1486), .CK(CLK), .RN(RST), .QN(n873) );
  DFFR_X1 \PC_TABLE_reg[12][18]  ( .D(n1467), .CK(CLK), .RN(RST), .QN(n854) );
  DFFR_X1 \PC_TABLE_reg[12][17]  ( .D(n1485), .CK(CLK), .RN(RST), .QN(n872) );
  DFFR_X1 \PC_TABLE_reg[12][16]  ( .D(n1468), .CK(CLK), .RN(RST), .QN(n855) );
  DFFR_X1 \PC_TABLE_reg[12][15]  ( .D(n1484), .CK(CLK), .RN(RST), .QN(n871) );
  DFFR_X1 \PC_TABLE_reg[12][13]  ( .D(n1483), .CK(CLK), .RN(RST), .QN(n870) );
  DFFR_X1 \PC_TABLE_reg[12][6]  ( .D(n1473), .CK(CLK), .RN(RST), .QN(n860) );
  DFFR_X1 \PC_TABLE_reg[12][0]  ( .D(n1476), .CK(CLK), .RN(RST), .QN(n863) );
  DFFR_X1 \PC_TABLE_reg[11][31]  ( .D(n1524), .CK(CLK), .RN(RST), .QN(n911) );
  DFFR_X1 \PC_TABLE_reg[11][28]  ( .D(n1494), .CK(CLK), .RN(RST), .QN(n881) );
  DFFR_X1 \PC_TABLE_reg[11][27]  ( .D(n1522), .CK(CLK), .RN(RST), .QN(n909) );
  DFFR_X1 \PC_TABLE_reg[11][22]  ( .D(n1497), .CK(CLK), .RN(RST), .QN(n884) );
  DFFR_X1 \PC_TABLE_reg[11][19]  ( .D(n1518), .CK(CLK), .RN(RST), .QN(n905) );
  DFFR_X1 \PC_TABLE_reg[11][17]  ( .D(n1517), .CK(CLK), .RN(RST), .QN(n904) );
  DFFR_X1 \PC_TABLE_reg[11][15]  ( .D(n1516), .CK(CLK), .RN(RST), .QN(n903) );
  DFFR_X1 \PC_TABLE_reg[11][12]  ( .D(n1502), .CK(CLK), .RN(RST), .QN(n889) );
  DFFR_X1 \PC_TABLE_reg[11][11]  ( .D(n1514), .CK(CLK), .RN(RST), .QN(n901) );
  DFFR_X1 \PC_TABLE_reg[11][8]  ( .D(n1504), .CK(CLK), .RN(RST), .QN(n891) );
  DFFR_X1 \PC_TABLE_reg[11][6]  ( .D(n1505), .CK(CLK), .RN(RST), .QN(n892) );
  DFFR_X1 \PC_TABLE_reg[11][0]  ( .D(n1508), .CK(CLK), .RN(RST), .QN(n895) );
  DFFR_X1 \PC_TABLE_reg[15][5]  ( .D(n1383), .CK(CLK), .RN(RST), .Q(n441), 
        .QN(n770) );
  DFFR_X1 \PC_TABLE_reg[15][4]  ( .D(n1379), .CK(CLK), .RN(RST), .Q(n425), 
        .QN(n766) );
  DFFR_X1 \PC_TABLE_reg[15][3]  ( .D(n1382), .CK(CLK), .RN(RST), .Q(n409), 
        .QN(n769) );
  DFFR_X1 \PC_TABLE_reg[15][2]  ( .D(n1380), .CK(CLK), .RN(RST), .Q(n393), 
        .QN(n767) );
  DFFR_X1 \PC_TABLE_reg[14][5]  ( .D(n1415), .CK(CLK), .RN(RST), .Q(n440), 
        .QN(n802) );
  DFFR_X1 \PC_TABLE_reg[14][4]  ( .D(n1410), .CK(CLK), .RN(RST), .Q(n424), 
        .QN(n797) );
  DFFR_X1 \PC_TABLE_reg[14][3]  ( .D(n1414), .CK(CLK), .RN(RST), .Q(n408), 
        .QN(n801) );
  DFFR_X1 \PC_TABLE_reg[7][18]  ( .D(n1627), .CK(CLK), .RN(RST), .QN(n1014) );
  DFFR_X1 \PC_TABLE_reg[7][26]  ( .D(n1623), .CK(CLK), .RN(RST), .QN(n1010) );
  DFFR_X1 \PC_TABLE_reg[7][24]  ( .D(n1624), .CK(CLK), .RN(RST), .QN(n1011) );
  DFFR_X1 \PC_TABLE_reg[7][22]  ( .D(n1625), .CK(CLK), .RN(RST), .QN(n1012) );
  DFFR_X1 \PC_TABLE_reg[10][28]  ( .D(n1526), .CK(CLK), .RN(RST), .QN(n913) );
  DFFR_X1 \PC_TABLE_reg[13][18]  ( .D(n1435), .CK(CLK), .RN(RST), .QN(n822) );
  DFFR_X1 \PC_TABLE_reg[11][18]  ( .D(n1499), .CK(CLK), .RN(RST), .QN(n886) );
  DFFR_X1 \PC_TABLE_reg[13][26]  ( .D(n1431), .CK(CLK), .RN(RST), .QN(n818) );
  DFFR_X1 \PC_TABLE_reg[10][26]  ( .D(n1527), .CK(CLK), .RN(RST), .QN(n914) );
  DFFR_X1 \PC_TABLE_reg[10][24]  ( .D(n1528), .CK(CLK), .RN(RST), .QN(n915) );
  DFFR_X1 \PC_TABLE_reg[10][22]  ( .D(n1529), .CK(CLK), .RN(RST), .QN(n916) );
  DFFR_X1 \PC_TABLE_reg[3][26]  ( .D(n1751), .CK(CLK), .RN(RST), .QN(n1138) );
  DFFR_X1 \PC_TABLE_reg[3][24]  ( .D(n1752), .CK(CLK), .RN(RST), .QN(n1139) );
  DFFR_X1 \PC_TABLE_reg[3][22]  ( .D(n1753), .CK(CLK), .RN(RST), .QN(n1140) );
  DFFR_X1 \PC_TABLE_reg[3][20]  ( .D(n1754), .CK(CLK), .RN(RST), .QN(n1141) );
  DFFR_X1 \PC_TABLE_reg[11][26]  ( .D(n1495), .CK(CLK), .RN(RST), .QN(n882) );
  DFFR_X1 \PC_TABLE_reg[13][24]  ( .D(n1432), .CK(CLK), .RN(RST), .QN(n819) );
  DFFR_X1 \PC_TABLE_reg[13][22]  ( .D(n1433), .CK(CLK), .RN(RST), .QN(n820) );
  DFFR_X1 \PC_TABLE_reg[11][24]  ( .D(n1496), .CK(CLK), .RN(RST), .QN(n883) );
  DFFR_X1 \PC_TABLE_reg[11][20]  ( .D(n1498), .CK(CLK), .RN(RST), .QN(n885) );
  DFFR_X1 \PC_TABLE_reg[10][27]  ( .D(n1554), .CK(CLK), .RN(RST), .QN(n941) );
  DFFR_X1 \PC_TABLE_reg[10][12]  ( .D(n1534), .CK(CLK), .RN(RST), .QN(n921) );
  DFFR_X1 \PC_TABLE_reg[10][11]  ( .D(n1546), .CK(CLK), .RN(RST), .QN(n933) );
  DFFR_X1 \PC_TABLE_reg[10][7]  ( .D(n1544), .CK(CLK), .RN(RST), .QN(n931) );
  DFFR_X1 \PC_TABLE_reg[10][1]  ( .D(n1541), .CK(CLK), .RN(RST), .QN(n928) );
  DFFR_X1 \PC_TABLE_reg[3][28]  ( .D(n1750), .CK(CLK), .RN(RST), .QN(n1137) );
  DFFR_X1 \PC_TABLE_reg[3][27]  ( .D(n1778), .CK(CLK), .RN(RST), .QN(n1165) );
  DFFR_X1 \PC_TABLE_reg[3][12]  ( .D(n1758), .CK(CLK), .RN(RST), .QN(n1145) );
  DFFR_X1 \PC_TABLE_reg[3][11]  ( .D(n1770), .CK(CLK), .RN(RST), .QN(n1157) );
  DFFR_X1 \PC_TABLE_reg[3][7]  ( .D(n1768), .CK(CLK), .RN(RST), .QN(n1155) );
  DFFR_X1 \PC_TABLE_reg[3][1]  ( .D(n1765), .CK(CLK), .RN(RST), .QN(n1152) );
  DFFR_X1 \PC_TABLE_reg[10][23]  ( .D(n1552), .CK(CLK), .RN(RST), .QN(n939) );
  DFFR_X1 \PC_TABLE_reg[10][21]  ( .D(n1551), .CK(CLK), .RN(RST), .QN(n938) );
  DFFR_X1 \PC_TABLE_reg[10][20]  ( .D(n1530), .CK(CLK), .RN(RST), .QN(n917) );
  DFFR_X1 \PC_TABLE_reg[10][19]  ( .D(n1550), .CK(CLK), .RN(RST), .QN(n937) );
  DFFR_X1 \PC_TABLE_reg[10][18]  ( .D(n1531), .CK(CLK), .RN(RST), .QN(n918) );
  DFFR_X1 \PC_TABLE_reg[10][17]  ( .D(n1549), .CK(CLK), .RN(RST), .QN(n936) );
  DFFR_X1 \PC_TABLE_reg[10][16]  ( .D(n1532), .CK(CLK), .RN(RST), .QN(n919) );
  DFFR_X1 \PC_TABLE_reg[10][15]  ( .D(n1548), .CK(CLK), .RN(RST), .QN(n935) );
  DFFR_X1 \PC_TABLE_reg[10][13]  ( .D(n1547), .CK(CLK), .RN(RST), .QN(n934) );
  DFFR_X1 \PC_TABLE_reg[10][6]  ( .D(n1537), .CK(CLK), .RN(RST), .QN(n924) );
  DFFR_X1 \PC_TABLE_reg[10][0]  ( .D(n1540), .CK(CLK), .RN(RST), .QN(n927) );
  DFFR_X1 \PC_TABLE_reg[3][23]  ( .D(n1776), .CK(CLK), .RN(RST), .QN(n1163) );
  DFFR_X1 \PC_TABLE_reg[3][21]  ( .D(n1775), .CK(CLK), .RN(RST), .QN(n1162) );
  DFFR_X1 \PC_TABLE_reg[3][19]  ( .D(n1774), .CK(CLK), .RN(RST), .QN(n1161) );
  DFFR_X1 \PC_TABLE_reg[3][18]  ( .D(n1755), .CK(CLK), .RN(RST), .QN(n1142) );
  DFFR_X1 \PC_TABLE_reg[3][17]  ( .D(n1773), .CK(CLK), .RN(RST), .QN(n1160) );
  DFFR_X1 \PC_TABLE_reg[3][16]  ( .D(n1756), .CK(CLK), .RN(RST), .QN(n1143) );
  DFFR_X1 \PC_TABLE_reg[3][15]  ( .D(n1772), .CK(CLK), .RN(RST), .QN(n1159) );
  DFFR_X1 \PC_TABLE_reg[3][13]  ( .D(n1771), .CK(CLK), .RN(RST), .QN(n1158) );
  DFFR_X1 \PC_TABLE_reg[3][6]  ( .D(n1761), .CK(CLK), .RN(RST), .QN(n1148) );
  DFFR_X1 \PC_TABLE_reg[3][0]  ( .D(n1764), .CK(CLK), .RN(RST), .QN(n1151) );
  DFFR_X1 \PC_TABLE_reg[10][31]  ( .D(n1556), .CK(CLK), .RN(RST), .QN(n943) );
  DFFR_X1 \PC_TABLE_reg[10][30]  ( .D(n1525), .CK(CLK), .RN(RST), .QN(n912) );
  DFFR_X1 \PC_TABLE_reg[10][29]  ( .D(n1555), .CK(CLK), .RN(RST), .QN(n942) );
  DFFR_X1 \PC_TABLE_reg[10][25]  ( .D(n1553), .CK(CLK), .RN(RST), .QN(n940) );
  DFFR_X1 \PC_TABLE_reg[10][14]  ( .D(n1533), .CK(CLK), .RN(RST), .QN(n920) );
  DFFR_X1 \PC_TABLE_reg[10][10]  ( .D(n1535), .CK(CLK), .RN(RST), .QN(n922) );
  DFFR_X1 \PC_TABLE_reg[10][9]  ( .D(n1545), .CK(CLK), .RN(RST), .QN(n932) );
  DFFR_X1 \PC_TABLE_reg[10][8]  ( .D(n1536), .CK(CLK), .RN(RST), .QN(n923) );
  DFFR_X1 \PC_TABLE_reg[3][31]  ( .D(n1780), .CK(CLK), .RN(RST), .QN(n1167) );
  DFFR_X1 \PC_TABLE_reg[3][30]  ( .D(n1749), .CK(CLK), .RN(RST), .QN(n1136) );
  DFFR_X1 \PC_TABLE_reg[3][29]  ( .D(n1779), .CK(CLK), .RN(RST), .QN(n1166) );
  DFFR_X1 \PC_TABLE_reg[3][25]  ( .D(n1777), .CK(CLK), .RN(RST), .QN(n1164) );
  DFFR_X1 \PC_TABLE_reg[3][14]  ( .D(n1757), .CK(CLK), .RN(RST), .QN(n1144) );
  DFFR_X1 \PC_TABLE_reg[3][10]  ( .D(n1759), .CK(CLK), .RN(RST), .QN(n1146) );
  DFFR_X1 \PC_TABLE_reg[3][9]  ( .D(n1769), .CK(CLK), .RN(RST), .QN(n1156) );
  DFFR_X1 \PC_TABLE_reg[3][8]  ( .D(n1760), .CK(CLK), .RN(RST), .QN(n1147) );
  DFFR_X1 \PC_TABLE_reg[15][20]  ( .D(n1371), .CK(CLK), .RN(RST), .Q(n681), 
        .QN(n758) );
  DFFR_X1 \PC_TABLE_reg[15][18]  ( .D(n1372), .CK(CLK), .RN(RST), .Q(n649), 
        .QN(n759) );
  DFFR_X1 \PC_TABLE_reg[15][26]  ( .D(n1368), .CK(CLK), .RN(RST), .Q(n265), 
        .QN(n755) );
  DFFR_X1 \PC_TABLE_reg[15][24]  ( .D(n1369), .CK(CLK), .RN(RST), .Q(n233), 
        .QN(n756) );
  DFFR_X1 \PC_TABLE_reg[14][0]  ( .D(n1412), .CK(CLK), .RN(RST), .Q(n360), 
        .QN(n799) );
  DFFR_X1 \PC_TABLE_reg[14][20]  ( .D(n1402), .CK(CLK), .RN(RST), .Q(n680), 
        .QN(n789) );
  DFFR_X1 \PC_TABLE_reg[14][26]  ( .D(n1399), .CK(CLK), .RN(RST), .Q(n264), 
        .QN(n786) );
  DFFR_X1 \PC_TABLE_reg[14][24]  ( .D(n1400), .CK(CLK), .RN(RST), .Q(n232), 
        .QN(n787) );
  DFFR_X1 \PC_TABLE_reg[15][0]  ( .D(n1877), .CK(CLK), .RN(RST), .Q(n361), 
        .QN(n1264) );
  DFFR_X1 \PC_TABLE_reg[15][31]  ( .D(n1396), .CK(CLK), .RN(RST), .Q(n345), 
        .QN(n783) );
  DFFR_X1 \PC_TABLE_reg[15][30]  ( .D(n1366), .CK(CLK), .RN(RST), .Q(n329), 
        .QN(n753) );
  DFFR_X1 \PC_TABLE_reg[15][29]  ( .D(n1395), .CK(CLK), .RN(RST), .Q(n313), 
        .QN(n782) );
  DFFR_X1 \PC_TABLE_reg[15][28]  ( .D(n1367), .CK(CLK), .RN(RST), .Q(n297), 
        .QN(n754) );
  DFFR_X1 \PC_TABLE_reg[15][27]  ( .D(n1394), .CK(CLK), .RN(RST), .Q(n281), 
        .QN(n781) );
  DFFR_X1 \PC_TABLE_reg[15][25]  ( .D(n1393), .CK(CLK), .RN(RST), .Q(n249), 
        .QN(n780) );
  DFFR_X1 \PC_TABLE_reg[15][23]  ( .D(n1392), .CK(CLK), .RN(RST), .Q(n217), 
        .QN(n779) );
  DFFR_X1 \PC_TABLE_reg[15][22]  ( .D(n1370), .CK(CLK), .RN(RST), .Q(n201), 
        .QN(n757) );
  DFFR_X1 \PC_TABLE_reg[15][21]  ( .D(n1391), .CK(CLK), .RN(RST), .Q(n704), 
        .QN(n778) );
  DFFR_X1 \PC_TABLE_reg[15][19]  ( .D(n1390), .CK(CLK), .RN(RST), .Q(n665), 
        .QN(n777) );
  DFFR_X1 \PC_TABLE_reg[15][17]  ( .D(n1389), .CK(CLK), .RN(RST), .Q(n633), 
        .QN(n776) );
  DFFR_X1 \PC_TABLE_reg[15][16]  ( .D(n1373), .CK(CLK), .RN(RST), .Q(n617), 
        .QN(n760) );
  DFFR_X1 \PC_TABLE_reg[15][15]  ( .D(n1388), .CK(CLK), .RN(RST), .Q(n601), 
        .QN(n775) );
  DFFR_X1 \PC_TABLE_reg[15][14]  ( .D(n1374), .CK(CLK), .RN(RST), .Q(n585), 
        .QN(n761) );
  DFFR_X1 \PC_TABLE_reg[15][13]  ( .D(n1387), .CK(CLK), .RN(RST), .Q(n569), 
        .QN(n774) );
  DFFR_X1 \PC_TABLE_reg[15][12]  ( .D(n1375), .CK(CLK), .RN(RST), .Q(n553), 
        .QN(n762) );
  DFFR_X1 \PC_TABLE_reg[15][11]  ( .D(n1386), .CK(CLK), .RN(RST), .Q(n537), 
        .QN(n773) );
  DFFR_X1 \PC_TABLE_reg[15][10]  ( .D(n1376), .CK(CLK), .RN(RST), .Q(n521), 
        .QN(n763) );
  DFFR_X1 \PC_TABLE_reg[15][9]  ( .D(n1385), .CK(CLK), .RN(RST), .Q(n505), 
        .QN(n772) );
  DFFR_X1 \PC_TABLE_reg[15][8]  ( .D(n1377), .CK(CLK), .RN(RST), .Q(n489), 
        .QN(n764) );
  DFFR_X1 \PC_TABLE_reg[15][7]  ( .D(n1384), .CK(CLK), .RN(RST), .Q(n473), 
        .QN(n771) );
  DFFR_X1 \PC_TABLE_reg[15][6]  ( .D(n1378), .CK(CLK), .RN(RST), .Q(n457), 
        .QN(n765) );
  DFFR_X1 \PC_TABLE_reg[15][1]  ( .D(n1381), .CK(CLK), .RN(RST), .Q(n377), 
        .QN(n768) );
  DFFR_X1 \PC_TABLE_reg[14][31]  ( .D(n1428), .CK(CLK), .RN(RST), .Q(n344), 
        .QN(n815) );
  DFFR_X1 \PC_TABLE_reg[14][30]  ( .D(n1397), .CK(CLK), .RN(RST), .Q(n328), 
        .QN(n784) );
  DFFR_X1 \PC_TABLE_reg[14][29]  ( .D(n1427), .CK(CLK), .RN(RST), .Q(n312), 
        .QN(n814) );
  DFFR_X1 \PC_TABLE_reg[14][27]  ( .D(n1426), .CK(CLK), .RN(RST), .Q(n280), 
        .QN(n813) );
  DFFR_X1 \PC_TABLE_reg[14][25]  ( .D(n1425), .CK(CLK), .RN(RST), .Q(n248), 
        .QN(n812) );
  DFFR_X1 \PC_TABLE_reg[14][23]  ( .D(n1424), .CK(CLK), .RN(RST), .Q(n216), 
        .QN(n811) );
  DFFR_X1 \PC_TABLE_reg[14][21]  ( .D(n1423), .CK(CLK), .RN(RST), .Q(n703), 
        .QN(n810) );
  DFFR_X1 \PC_TABLE_reg[14][19]  ( .D(n1422), .CK(CLK), .RN(RST), .Q(n664), 
        .QN(n809) );
  DFFR_X1 \PC_TABLE_reg[14][18]  ( .D(n1403), .CK(CLK), .RN(RST), .Q(n648), 
        .QN(n790) );
  DFFR_X1 \PC_TABLE_reg[14][17]  ( .D(n1421), .CK(CLK), .RN(RST), .Q(n632), 
        .QN(n808) );
  DFFR_X1 \PC_TABLE_reg[14][16]  ( .D(n1404), .CK(CLK), .RN(RST), .Q(n616), 
        .QN(n791) );
  DFFR_X1 \PC_TABLE_reg[14][15]  ( .D(n1420), .CK(CLK), .RN(RST), .Q(n600), 
        .QN(n807) );
  DFFR_X1 \PC_TABLE_reg[14][14]  ( .D(n1405), .CK(CLK), .RN(RST), .Q(n584), 
        .QN(n792) );
  DFFR_X1 \PC_TABLE_reg[14][13]  ( .D(n1419), .CK(CLK), .RN(RST), .Q(n568), 
        .QN(n806) );
  DFFR_X1 \PC_TABLE_reg[14][12]  ( .D(n1406), .CK(CLK), .RN(RST), .Q(n552), 
        .QN(n793) );
  DFFR_X1 \PC_TABLE_reg[14][11]  ( .D(n1418), .CK(CLK), .RN(RST), .Q(n536), 
        .QN(n805) );
  DFFR_X1 \PC_TABLE_reg[14][10]  ( .D(n1407), .CK(CLK), .RN(RST), .Q(n520), 
        .QN(n794) );
  DFFR_X1 \PC_TABLE_reg[14][9]  ( .D(n1417), .CK(CLK), .RN(RST), .Q(n504), 
        .QN(n804) );
  DFFR_X1 \PC_TABLE_reg[14][8]  ( .D(n1408), .CK(CLK), .RN(RST), .Q(n488), 
        .QN(n795) );
  DFFR_X1 \PC_TABLE_reg[14][7]  ( .D(n1416), .CK(CLK), .RN(RST), .Q(n472), 
        .QN(n803) );
  DFFR_X1 \PC_TABLE_reg[14][6]  ( .D(n1409), .CK(CLK), .RN(RST), .Q(n456), 
        .QN(n796) );
  DFFR_X1 \PC_TABLE_reg[14][1]  ( .D(n1413), .CK(CLK), .RN(RST), .Q(n376), 
        .QN(n800) );
  DFFR_X1 \PC_TABLE_reg[14][28]  ( .D(n1398), .CK(CLK), .RN(RST), .Q(n296), 
        .QN(n785) );
  DFFR_X1 \PC_TABLE_reg[14][22]  ( .D(n1401), .CK(CLK), .RN(RST), .Q(n200), 
        .QN(n788) );
  DFFR_X1 \PC_TABLE_reg[9][28]  ( .D(n1558), .CK(CLK), .RN(RST), .Q(n300), 
        .QN(n945) );
  DFFR_X1 \PC_TABLE_reg[9][26]  ( .D(n1559), .CK(CLK), .RN(RST), .Q(n268), 
        .QN(n946) );
  DFFR_X1 \PC_TABLE_reg[9][24]  ( .D(n1560), .CK(CLK), .RN(RST), .Q(n236), 
        .QN(n947) );
  DFFR_X1 \PC_TABLE_reg[9][22]  ( .D(n1561), .CK(CLK), .RN(RST), .Q(n204), 
        .QN(n948) );
  DFFR_X1 \PC_TABLE_reg[9][20]  ( .D(n1562), .CK(CLK), .RN(RST), .Q(n684), 
        .QN(n949) );
  DFFR_X1 \PC_TABLE_reg[9][18]  ( .D(n1563), .CK(CLK), .RN(RST), .Q(n652), 
        .QN(n950) );
  DFFR_X1 \PC_TABLE_reg[5][28]  ( .D(n1686), .CK(CLK), .RN(RST), .Q(n291), 
        .QN(n1073) );
  DFFR_X1 \PC_TABLE_reg[5][26]  ( .D(n1687), .CK(CLK), .RN(RST), .Q(n259), 
        .QN(n1074) );
  DFFR_X1 \PC_TABLE_reg[5][24]  ( .D(n1688), .CK(CLK), .RN(RST), .Q(n227), 
        .QN(n1075) );
  DFFR_X1 \PC_TABLE_reg[5][22]  ( .D(n1689), .CK(CLK), .RN(RST), .Q(n195), 
        .QN(n1076) );
  DFFR_X1 \PC_TABLE_reg[5][20]  ( .D(n1690), .CK(CLK), .RN(RST), .Q(n675), 
        .QN(n1077) );
  DFFR_X1 \PC_TABLE_reg[5][18]  ( .D(n1691), .CK(CLK), .RN(RST), .Q(n643), 
        .QN(n1078) );
  DFFR_X1 \PC_TABLE_reg[8][28]  ( .D(n1590), .CK(CLK), .RN(RST), .Q(n299), 
        .QN(n977) );
  DFFR_X1 \PC_TABLE_reg[8][26]  ( .D(n1591), .CK(CLK), .RN(RST), .Q(n267), 
        .QN(n978) );
  DFFR_X1 \PC_TABLE_reg[8][24]  ( .D(n1592), .CK(CLK), .RN(RST), .Q(n235), 
        .QN(n979) );
  DFFR_X1 \PC_TABLE_reg[8][22]  ( .D(n1593), .CK(CLK), .RN(RST), .Q(n203), 
        .QN(n980) );
  DFFR_X1 \PC_TABLE_reg[8][20]  ( .D(n1594), .CK(CLK), .RN(RST), .Q(n683), 
        .QN(n981) );
  DFFR_X1 \PC_TABLE_reg[8][18]  ( .D(n1595), .CK(CLK), .RN(RST), .Q(n651), 
        .QN(n982) );
  DFFR_X1 \PC_TABLE_reg[8][16]  ( .D(n1596), .CK(CLK), .RN(RST), .Q(n619), 
        .QN(n983) );
  DFFR_X1 \PC_TABLE_reg[4][28]  ( .D(n1718), .CK(CLK), .RN(RST), .Q(n290), 
        .QN(n1105) );
  DFFR_X1 \PC_TABLE_reg[4][26]  ( .D(n1719), .CK(CLK), .RN(RST), .Q(n258), 
        .QN(n1106) );
  DFFR_X1 \PC_TABLE_reg[4][24]  ( .D(n1720), .CK(CLK), .RN(RST), .Q(n226), 
        .QN(n1107) );
  DFFR_X1 \PC_TABLE_reg[4][22]  ( .D(n1721), .CK(CLK), .RN(RST), .Q(n194), 
        .QN(n1108) );
  DFFR_X1 \PC_TABLE_reg[4][20]  ( .D(n1722), .CK(CLK), .RN(RST), .Q(n674), 
        .QN(n1109) );
  DFFR_X1 \PC_TABLE_reg[4][18]  ( .D(n1723), .CK(CLK), .RN(RST), .Q(n642), 
        .QN(n1110) );
  DFFR_X1 \PC_TABLE_reg[4][16]  ( .D(n1724), .CK(CLK), .RN(RST), .Q(n610), 
        .QN(n1111) );
  DFFR_X1 \PC_TABLE_reg[1][28]  ( .D(n1814), .CK(CLK), .RN(RST), .Q(n294), 
        .QN(n1201) );
  DFFR_X1 \PC_TABLE_reg[1][26]  ( .D(n1815), .CK(CLK), .RN(RST), .Q(n262), 
        .QN(n1202) );
  DFFR_X1 \PC_TABLE_reg[1][24]  ( .D(n1816), .CK(CLK), .RN(RST), .Q(n230), 
        .QN(n1203) );
  DFFR_X1 \PC_TABLE_reg[1][22]  ( .D(n1817), .CK(CLK), .RN(RST), .Q(n198), 
        .QN(n1204) );
  DFFR_X1 \PC_TABLE_reg[1][20]  ( .D(n1818), .CK(CLK), .RN(RST), .Q(n678), 
        .QN(n1205) );
  DFFR_X1 \PC_TABLE_reg[1][18]  ( .D(n1819), .CK(CLK), .RN(RST), .Q(n646), 
        .QN(n1206) );
  DFFR_X1 \PC_TABLE_reg[1][16]  ( .D(n1820), .CK(CLK), .RN(RST), .Q(n614), 
        .QN(n1207) );
  DFFR_X1 \PC_TABLE_reg[8][30]  ( .D(n1589), .CK(CLK), .RN(RST), .Q(n331), 
        .QN(n976) );
  DFFR_X1 \PC_TABLE_reg[8][29]  ( .D(n1619), .CK(CLK), .RN(RST), .Q(n315), 
        .QN(n1006) );
  DFFR_X1 \PC_TABLE_reg[8][27]  ( .D(n1618), .CK(CLK), .RN(RST), .Q(n283), 
        .QN(n1005) );
  DFFR_X1 \PC_TABLE_reg[8][23]  ( .D(n1616), .CK(CLK), .RN(RST), .Q(n219), 
        .QN(n1003) );
  DFFR_X1 \PC_TABLE_reg[8][21]  ( .D(n1615), .CK(CLK), .RN(RST), .Q(n708), 
        .QN(n1002) );
  DFFR_X1 \PC_TABLE_reg[8][19]  ( .D(n1614), .CK(CLK), .RN(RST), .Q(n667), 
        .QN(n1001) );
  DFFR_X1 \PC_TABLE_reg[8][17]  ( .D(n1613), .CK(CLK), .RN(RST), .Q(n635), 
        .QN(n1000) );
  DFFR_X1 \PC_TABLE_reg[8][15]  ( .D(n1612), .CK(CLK), .RN(RST), .Q(n603), 
        .QN(n999) );
  DFFR_X1 \PC_TABLE_reg[8][11]  ( .D(n1610), .CK(CLK), .RN(RST), .Q(n539), 
        .QN(n997) );
  DFFR_X1 \PC_TABLE_reg[4][30]  ( .D(n1717), .CK(CLK), .RN(RST), .Q(n322), 
        .QN(n1104) );
  DFFR_X1 \PC_TABLE_reg[4][29]  ( .D(n1747), .CK(CLK), .RN(RST), .Q(n306), 
        .QN(n1134) );
  DFFR_X1 \PC_TABLE_reg[4][27]  ( .D(n1746), .CK(CLK), .RN(RST), .Q(n274), 
        .QN(n1133) );
  DFFR_X1 \PC_TABLE_reg[4][23]  ( .D(n1744), .CK(CLK), .RN(RST), .Q(n210), 
        .QN(n1131) );
  DFFR_X1 \PC_TABLE_reg[4][21]  ( .D(n1743), .CK(CLK), .RN(RST), .Q(n690), 
        .QN(n1130) );
  DFFR_X1 \PC_TABLE_reg[4][19]  ( .D(n1742), .CK(CLK), .RN(RST), .Q(n658), 
        .QN(n1129) );
  DFFR_X1 \PC_TABLE_reg[4][17]  ( .D(n1741), .CK(CLK), .RN(RST), .Q(n626), 
        .QN(n1128) );
  DFFR_X1 \PC_TABLE_reg[4][15]  ( .D(n1740), .CK(CLK), .RN(RST), .Q(n594), 
        .QN(n1127) );
  DFFR_X1 \PC_TABLE_reg[4][11]  ( .D(n1738), .CK(CLK), .RN(RST), .Q(n530), 
        .QN(n1125) );
  DFFR_X1 \PC_TABLE_reg[1][30]  ( .D(n1813), .CK(CLK), .RN(RST), .Q(n326), 
        .QN(n1200) );
  DFFR_X1 \PC_TABLE_reg[1][29]  ( .D(n1843), .CK(CLK), .RN(RST), .Q(n310), 
        .QN(n1230) );
  DFFR_X1 \PC_TABLE_reg[1][27]  ( .D(n1842), .CK(CLK), .RN(RST), .Q(n278), 
        .QN(n1229) );
  DFFR_X1 \PC_TABLE_reg[1][23]  ( .D(n1840), .CK(CLK), .RN(RST), .Q(n214), 
        .QN(n1227) );
  DFFR_X1 \PC_TABLE_reg[1][21]  ( .D(n1839), .CK(CLK), .RN(RST), .Q(n700), 
        .QN(n1226) );
  DFFR_X1 \PC_TABLE_reg[1][19]  ( .D(n1838), .CK(CLK), .RN(RST), .Q(n662), 
        .QN(n1225) );
  DFFR_X1 \PC_TABLE_reg[1][17]  ( .D(n1837), .CK(CLK), .RN(RST), .Q(n630), 
        .QN(n1224) );
  DFFR_X1 \PC_TABLE_reg[1][15]  ( .D(n1836), .CK(CLK), .RN(RST), .Q(n598), 
        .QN(n1223) );
  DFFR_X1 \PC_TABLE_reg[1][11]  ( .D(n1834), .CK(CLK), .RN(RST), .Q(n534), 
        .QN(n1221) );
  DFFR_X1 \PC_TABLE_reg[8][0]  ( .D(n1604), .CK(CLK), .RN(RST), .Q(n363), .QN(
        n991) );
  DFFR_X1 \PC_TABLE_reg[4][0]  ( .D(n1732), .CK(CLK), .RN(RST), .Q(n354), .QN(
        n1119) );
  DFFR_X1 \PC_TABLE_reg[8][31]  ( .D(n1620), .CK(CLK), .RN(RST), .Q(n347), 
        .QN(n1007) );
  DFFR_X1 \PC_TABLE_reg[8][25]  ( .D(n1617), .CK(CLK), .RN(RST), .Q(n251), 
        .QN(n1004) );
  DFFR_X1 \PC_TABLE_reg[8][14]  ( .D(n1597), .CK(CLK), .RN(RST), .Q(n587), 
        .QN(n984) );
  DFFR_X1 \PC_TABLE_reg[8][13]  ( .D(n1611), .CK(CLK), .RN(RST), .Q(n571), 
        .QN(n998) );
  DFFR_X1 \PC_TABLE_reg[8][12]  ( .D(n1598), .CK(CLK), .RN(RST), .Q(n555), 
        .QN(n985) );
  DFFR_X1 \PC_TABLE_reg[8][10]  ( .D(n1599), .CK(CLK), .RN(RST), .Q(n523), 
        .QN(n986) );
  DFFR_X1 \PC_TABLE_reg[8][9]  ( .D(n1609), .CK(CLK), .RN(RST), .Q(n507), .QN(
        n996) );
  DFFR_X1 \PC_TABLE_reg[8][8]  ( .D(n1600), .CK(CLK), .RN(RST), .Q(n491), .QN(
        n987) );
  DFFR_X1 \PC_TABLE_reg[8][7]  ( .D(n1608), .CK(CLK), .RN(RST), .Q(n475), .QN(
        n995) );
  DFFR_X1 \PC_TABLE_reg[8][6]  ( .D(n1601), .CK(CLK), .RN(RST), .Q(n459), .QN(
        n988) );
  DFFR_X1 \PC_TABLE_reg[4][31]  ( .D(n1748), .CK(CLK), .RN(RST), .Q(n338), 
        .QN(n1135) );
  DFFR_X1 \PC_TABLE_reg[4][25]  ( .D(n1745), .CK(CLK), .RN(RST), .Q(n242), 
        .QN(n1132) );
  DFFR_X1 \PC_TABLE_reg[4][14]  ( .D(n1725), .CK(CLK), .RN(RST), .Q(n578), 
        .QN(n1112) );
  DFFR_X1 \PC_TABLE_reg[4][13]  ( .D(n1739), .CK(CLK), .RN(RST), .Q(n562), 
        .QN(n1126) );
  DFFR_X1 \PC_TABLE_reg[4][12]  ( .D(n1726), .CK(CLK), .RN(RST), .Q(n546), 
        .QN(n1113) );
  DFFR_X1 \PC_TABLE_reg[4][10]  ( .D(n1727), .CK(CLK), .RN(RST), .Q(n514), 
        .QN(n1114) );
  DFFR_X1 \PC_TABLE_reg[4][9]  ( .D(n1737), .CK(CLK), .RN(RST), .Q(n498), .QN(
        n1124) );
  DFFR_X1 \PC_TABLE_reg[4][8]  ( .D(n1728), .CK(CLK), .RN(RST), .Q(n482), .QN(
        n1115) );
  DFFR_X1 \PC_TABLE_reg[4][7]  ( .D(n1736), .CK(CLK), .RN(RST), .Q(n466), .QN(
        n1123) );
  DFFR_X1 \PC_TABLE_reg[4][6]  ( .D(n1729), .CK(CLK), .RN(RST), .Q(n450), .QN(
        n1116) );
  DFFR_X1 \PC_TABLE_reg[8][1]  ( .D(n1605), .CK(CLK), .RN(RST), .Q(n379), .QN(
        n992) );
  DFFR_X1 \PC_TABLE_reg[4][1]  ( .D(n1733), .CK(CLK), .RN(RST), .Q(n370), .QN(
        n1120) );
  DFFR_X1 \PC_TABLE_reg[1][0]  ( .D(n1828), .CK(CLK), .RN(RST), .Q(n358), .QN(
        n1215) );
  DFFR_X1 \PC_TABLE_reg[1][31]  ( .D(n1844), .CK(CLK), .RN(RST), .Q(n342), 
        .QN(n1231) );
  DFFR_X1 \PC_TABLE_reg[1][25]  ( .D(n1841), .CK(CLK), .RN(RST), .Q(n246), 
        .QN(n1228) );
  DFFR_X1 \PC_TABLE_reg[1][14]  ( .D(n1821), .CK(CLK), .RN(RST), .Q(n582), 
        .QN(n1208) );
  DFFR_X1 \PC_TABLE_reg[1][13]  ( .D(n1835), .CK(CLK), .RN(RST), .Q(n566), 
        .QN(n1222) );
  DFFR_X1 \PC_TABLE_reg[1][12]  ( .D(n1822), .CK(CLK), .RN(RST), .Q(n550), 
        .QN(n1209) );
  DFFR_X1 \PC_TABLE_reg[1][10]  ( .D(n1823), .CK(CLK), .RN(RST), .Q(n518), 
        .QN(n1210) );
  DFFR_X1 \PC_TABLE_reg[1][9]  ( .D(n1833), .CK(CLK), .RN(RST), .Q(n502), .QN(
        n1220) );
  DFFR_X1 \PC_TABLE_reg[1][8]  ( .D(n1824), .CK(CLK), .RN(RST), .Q(n486), .QN(
        n1211) );
  DFFR_X1 \PC_TABLE_reg[1][7]  ( .D(n1832), .CK(CLK), .RN(RST), .Q(n470), .QN(
        n1219) );
  DFFR_X1 \PC_TABLE_reg[1][6]  ( .D(n1825), .CK(CLK), .RN(RST), .Q(n454), .QN(
        n1212) );
  DFFR_X1 \PC_TABLE_reg[1][1]  ( .D(n1829), .CK(CLK), .RN(RST), .Q(n374), .QN(
        n1216) );
  DFFR_X1 \PC_TABLE_reg[9][0]  ( .D(n1572), .CK(CLK), .RN(RST), .Q(n364), .QN(
        n959) );
  DFFR_X1 \PC_TABLE_reg[5][0]  ( .D(n1700), .CK(CLK), .RN(RST), .Q(n355), .QN(
        n1087) );
  DFFR_X1 \PC_TABLE_reg[9][31]  ( .D(n1588), .CK(CLK), .RN(RST), .Q(n348), 
        .QN(n975) );
  DFFR_X1 \PC_TABLE_reg[9][16]  ( .D(n1564), .CK(CLK), .RN(RST), .Q(n620), 
        .QN(n951) );
  DFFR_X1 \PC_TABLE_reg[9][15]  ( .D(n1580), .CK(CLK), .RN(RST), .Q(n604), 
        .QN(n967) );
  DFFR_X1 \PC_TABLE_reg[9][14]  ( .D(n1565), .CK(CLK), .RN(RST), .Q(n588), 
        .QN(n952) );
  DFFR_X1 \PC_TABLE_reg[9][12]  ( .D(n1566), .CK(CLK), .RN(RST), .Q(n556), 
        .QN(n953) );
  DFFR_X1 \PC_TABLE_reg[9][10]  ( .D(n1567), .CK(CLK), .RN(RST), .Q(n524), 
        .QN(n954) );
  DFFR_X1 \PC_TABLE_reg[9][9]  ( .D(n1577), .CK(CLK), .RN(RST), .Q(n508), .QN(
        n964) );
  DFFR_X1 \PC_TABLE_reg[9][8]  ( .D(n1568), .CK(CLK), .RN(RST), .Q(n492), .QN(
        n955) );
  DFFR_X1 \PC_TABLE_reg[9][7]  ( .D(n1576), .CK(CLK), .RN(RST), .Q(n476), .QN(
        n963) );
  DFFR_X1 \PC_TABLE_reg[9][6]  ( .D(n1569), .CK(CLK), .RN(RST), .Q(n460), .QN(
        n956) );
  DFFR_X1 \PC_TABLE_reg[5][31]  ( .D(n1716), .CK(CLK), .RN(RST), .Q(n339), 
        .QN(n1103) );
  DFFR_X1 \PC_TABLE_reg[5][16]  ( .D(n1692), .CK(CLK), .RN(RST), .Q(n611), 
        .QN(n1079) );
  DFFR_X1 \PC_TABLE_reg[5][15]  ( .D(n1708), .CK(CLK), .RN(RST), .Q(n595), 
        .QN(n1095) );
  DFFR_X1 \PC_TABLE_reg[5][14]  ( .D(n1693), .CK(CLK), .RN(RST), .Q(n579), 
        .QN(n1080) );
  DFFR_X1 \PC_TABLE_reg[5][12]  ( .D(n1694), .CK(CLK), .RN(RST), .Q(n547), 
        .QN(n1081) );
  DFFR_X1 \PC_TABLE_reg[5][10]  ( .D(n1695), .CK(CLK), .RN(RST), .Q(n515), 
        .QN(n1082) );
  DFFR_X1 \PC_TABLE_reg[5][9]  ( .D(n1705), .CK(CLK), .RN(RST), .Q(n499), .QN(
        n1092) );
  DFFR_X1 \PC_TABLE_reg[5][8]  ( .D(n1696), .CK(CLK), .RN(RST), .Q(n483), .QN(
        n1083) );
  DFFR_X1 \PC_TABLE_reg[5][7]  ( .D(n1704), .CK(CLK), .RN(RST), .Q(n467), .QN(
        n1091) );
  DFFR_X1 \PC_TABLE_reg[5][6]  ( .D(n1697), .CK(CLK), .RN(RST), .Q(n451), .QN(
        n1084) );
  DFFR_X1 \PC_TABLE_reg[9][1]  ( .D(n1573), .CK(CLK), .RN(RST), .Q(n380), .QN(
        n960) );
  DFFR_X1 \PC_TABLE_reg[5][1]  ( .D(n1701), .CK(CLK), .RN(RST), .Q(n371), .QN(
        n1088) );
  DFFR_X1 \PC_TABLE_reg[0][30]  ( .D(n1845), .CK(CLK), .RN(RST), .Q(n325), 
        .QN(n1232) );
  DFFR_X1 \PC_TABLE_reg[0][29]  ( .D(n1875), .CK(CLK), .RN(RST), .Q(n309), 
        .QN(n1262) );
  DFFR_X1 \PC_TABLE_reg[0][28]  ( .D(n1846), .CK(CLK), .RN(RST), .Q(n293), 
        .QN(n1233) );
  DFFR_X1 \PC_TABLE_reg[0][27]  ( .D(n1874), .CK(CLK), .RN(RST), .Q(n277), 
        .QN(n1261) );
  DFFR_X1 \PC_TABLE_reg[0][26]  ( .D(n1847), .CK(CLK), .RN(RST), .Q(n261), 
        .QN(n1234) );
  DFFR_X1 \PC_TABLE_reg[0][25]  ( .D(n1873), .CK(CLK), .RN(RST), .Q(n245), 
        .QN(n1260) );
  DFFR_X1 \PC_TABLE_reg[0][24]  ( .D(n1848), .CK(CLK), .RN(RST), .Q(n229), 
        .QN(n1235) );
  DFFR_X1 \PC_TABLE_reg[0][23]  ( .D(n1872), .CK(CLK), .RN(RST), .Q(n213), 
        .QN(n1259) );
  DFFR_X1 \PC_TABLE_reg[0][22]  ( .D(n1849), .CK(CLK), .RN(RST), .Q(n197), 
        .QN(n1236) );
  DFFR_X1 \PC_TABLE_reg[0][21]  ( .D(n1871), .CK(CLK), .RN(RST), .Q(n699), 
        .QN(n1258) );
  DFFR_X1 \PC_TABLE_reg[0][20]  ( .D(n1850), .CK(CLK), .RN(RST), .Q(n677), 
        .QN(n1237) );
  DFFR_X1 \PC_TABLE_reg[0][19]  ( .D(n1870), .CK(CLK), .RN(RST), .Q(n661), 
        .QN(n1257) );
  DFFR_X1 \PC_TABLE_reg[0][18]  ( .D(n1851), .CK(CLK), .RN(RST), .Q(n645), 
        .QN(n1238) );
  DFFR_X1 \PC_TABLE_reg[0][16]  ( .D(n1852), .CK(CLK), .RN(RST), .Q(n613), 
        .QN(n1239) );
  DFFR_X1 \PC_TABLE_reg[0][15]  ( .D(n1868), .CK(CLK), .RN(RST), .Q(n597), 
        .QN(n1255) );
  DFFR_X1 \PC_TABLE_reg[0][14]  ( .D(n1853), .CK(CLK), .RN(RST), .Q(n581), 
        .QN(n1240) );
  DFFR_X1 \PC_TABLE_reg[9][30]  ( .D(n1557), .CK(CLK), .RN(RST), .Q(n332), 
        .QN(n944) );
  DFFR_X1 \PC_TABLE_reg[9][29]  ( .D(n1587), .CK(CLK), .RN(RST), .Q(n316), 
        .QN(n974) );
  DFFR_X1 \PC_TABLE_reg[9][27]  ( .D(n1586), .CK(CLK), .RN(RST), .Q(n284), 
        .QN(n973) );
  DFFR_X1 \PC_TABLE_reg[9][25]  ( .D(n1585), .CK(CLK), .RN(RST), .Q(n252), 
        .QN(n972) );
  DFFR_X1 \PC_TABLE_reg[9][23]  ( .D(n1584), .CK(CLK), .RN(RST), .Q(n220), 
        .QN(n971) );
  DFFR_X1 \PC_TABLE_reg[9][21]  ( .D(n1583), .CK(CLK), .RN(RST), .Q(n709), 
        .QN(n970) );
  DFFR_X1 \PC_TABLE_reg[9][19]  ( .D(n1582), .CK(CLK), .RN(RST), .Q(n668), 
        .QN(n969) );
  DFFR_X1 \PC_TABLE_reg[9][17]  ( .D(n1581), .CK(CLK), .RN(RST), .Q(n636), 
        .QN(n968) );
  DFFR_X1 \PC_TABLE_reg[9][13]  ( .D(n1579), .CK(CLK), .RN(RST), .Q(n572), 
        .QN(n966) );
  DFFR_X1 \PC_TABLE_reg[9][11]  ( .D(n1578), .CK(CLK), .RN(RST), .Q(n540), 
        .QN(n965) );
  DFFR_X1 \PC_TABLE_reg[5][30]  ( .D(n1685), .CK(CLK), .RN(RST), .Q(n323), 
        .QN(n1072) );
  DFFR_X1 \PC_TABLE_reg[5][29]  ( .D(n1715), .CK(CLK), .RN(RST), .Q(n307), 
        .QN(n1102) );
  DFFR_X1 \PC_TABLE_reg[5][27]  ( .D(n1714), .CK(CLK), .RN(RST), .Q(n275), 
        .QN(n1101) );
  DFFR_X1 \PC_TABLE_reg[5][25]  ( .D(n1713), .CK(CLK), .RN(RST), .Q(n243), 
        .QN(n1100) );
  DFFR_X1 \PC_TABLE_reg[5][23]  ( .D(n1712), .CK(CLK), .RN(RST), .Q(n211), 
        .QN(n1099) );
  DFFR_X1 \PC_TABLE_reg[5][21]  ( .D(n1711), .CK(CLK), .RN(RST), .Q(n691), 
        .QN(n1098) );
  DFFR_X1 \PC_TABLE_reg[5][19]  ( .D(n1710), .CK(CLK), .RN(RST), .Q(n659), 
        .QN(n1097) );
  DFFR_X1 \PC_TABLE_reg[5][17]  ( .D(n1709), .CK(CLK), .RN(RST), .Q(n627), 
        .QN(n1096) );
  DFFR_X1 \PC_TABLE_reg[5][13]  ( .D(n1707), .CK(CLK), .RN(RST), .Q(n563), 
        .QN(n1094) );
  DFFR_X1 \PC_TABLE_reg[5][11]  ( .D(n1706), .CK(CLK), .RN(RST), .Q(n531), 
        .QN(n1093) );
  DFFR_X1 \PC_TABLE_reg[0][0]  ( .D(n1860), .CK(CLK), .RN(RST), .Q(n357), .QN(
        n1247) );
  DFFR_X1 \PC_TABLE_reg[0][31]  ( .D(n1876), .CK(CLK), .RN(RST), .Q(n341), 
        .QN(n1263) );
  DFFR_X1 \PC_TABLE_reg[0][17]  ( .D(n1869), .CK(CLK), .RN(RST), .Q(n629), 
        .QN(n1256) );
  DFFR_X1 \PC_TABLE_reg[0][13]  ( .D(n1867), .CK(CLK), .RN(RST), .Q(n565), 
        .QN(n1254) );
  DFFR_X1 \PC_TABLE_reg[0][12]  ( .D(n1854), .CK(CLK), .RN(RST), .Q(n549), 
        .QN(n1241) );
  DFFR_X1 \PC_TABLE_reg[0][11]  ( .D(n1866), .CK(CLK), .RN(RST), .Q(n533), 
        .QN(n1253) );
  DFFR_X1 \PC_TABLE_reg[0][10]  ( .D(n1855), .CK(CLK), .RN(RST), .Q(n517), 
        .QN(n1242) );
  DFFR_X1 \PC_TABLE_reg[0][9]  ( .D(n1865), .CK(CLK), .RN(RST), .Q(n501), .QN(
        n1252) );
  DFFR_X1 \PC_TABLE_reg[0][8]  ( .D(n1856), .CK(CLK), .RN(RST), .Q(n485), .QN(
        n1243) );
  DFFR_X1 \PC_TABLE_reg[0][7]  ( .D(n1864), .CK(CLK), .RN(RST), .Q(n469), .QN(
        n1251) );
  DFFR_X1 \PC_TABLE_reg[0][6]  ( .D(n1857), .CK(CLK), .RN(RST), .Q(n453), .QN(
        n1244) );
  DFFR_X1 \PC_TABLE_reg[0][1]  ( .D(n1861), .CK(CLK), .RN(RST), .Q(n373), .QN(
        n1248) );
  DFFR_X1 \PRED_HISTORY_reg[1][32]  ( .D(\PRED_HISTORY[0][32] ), .CK(CLK), 
        .RN(RST), .Q(MISS_HIT[1]), .QN(n749) );
  DFFR_X1 \PC_HISTORY_reg[1][3]  ( .D(\PC_HISTORY[0][3] ), .CK(CLK), .RN(RST), 
        .Q(\PC_HISTORY[1][3] ), .QN(n750) );
  DFFR_X1 \PC_HISTORY_reg[1][2]  ( .D(\PC_HISTORY[0][2] ), .CK(CLK), .RN(RST), 
        .Q(\PC_HISTORY[1][2] ), .QN(n748) );
  DFFR_X1 \PC_HISTORY_reg[1][1]  ( .D(\PC_HISTORY[0][1] ), .CK(CLK), .RN(RST), 
        .Q(\PC_HISTORY[1][1] ), .QN(n747) );
  DFFR_X1 \PC_HISTORY_reg[1][0]  ( .D(\PC_HISTORY[0][0] ), .CK(CLK), .RN(RST), 
        .Q(\PC_HISTORY[1][0] ), .QN(n751) );
  DFFR_X1 \PRED_TABLE_reg[15][1]  ( .D(n1360), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[15][1] ), .QN(n752) );
  DFFR_X1 \PRED_TABLE_reg[14][1]  ( .D(n1288), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[14][1] ), .QN(n739) );
  DFFR_X1 \PRED_TABLE_reg[13][1]  ( .D(n1287), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[13][1] ), .QN(n738) );
  DFFR_X1 \PRED_TABLE_reg[12][1]  ( .D(n1289), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[12][1] ), .QN(n740) );
  DFFR_X1 \PRED_TABLE_reg[11][1]  ( .D(n1286), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[11][1] ), .QN(n737) );
  DFFR_X1 \PRED_TABLE_reg[10][1]  ( .D(n1290), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[10][1] ), .QN(n741) );
  DFFR_X1 \PRED_TABLE_reg[9][1]  ( .D(n1285), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[9][1] ), .QN(n736) );
  DFFR_X1 \PRED_TABLE_reg[8][1]  ( .D(n1291), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[8][1] ), .QN(n742) );
  DFFR_X1 \PRED_TABLE_reg[7][1]  ( .D(n1284), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[7][1] ), .QN(n735) );
  DFFR_X1 \PRED_TABLE_reg[6][1]  ( .D(n1292), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[6][1] ), .QN(n743) );
  DFFR_X1 \PRED_TABLE_reg[5][1]  ( .D(n1283), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[5][1] ), .QN(n734) );
  DFFR_X1 \PRED_TABLE_reg[4][1]  ( .D(n1293), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[4][1] ), .QN(n744) );
  DFFR_X1 \PRED_TABLE_reg[3][1]  ( .D(n1282), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[3][1] ), .QN(n733) );
  DFFR_X1 \PRED_TABLE_reg[2][1]  ( .D(n1294), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[2][1] ), .QN(n745) );
  DFFR_X1 \PRED_TABLE_reg[1][1]  ( .D(n1281), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[1][1] ), .QN(n732) );
  DFFR_X1 \PRED_TABLE_reg[0][1]  ( .D(n1295), .CK(CLK), .RN(RST), .Q(
        \PRED_TABLE[0][1] ), .QN(n746) );
  DFFR_X2 \PRED_HISTORY_reg[0][31]  ( .D(PRED[31]), .CK(CLK), .RN(n2207), .Q(
        \PRED_HISTORY[0][31] ) );
  INV_X1 U3 ( .A(n404), .ZN(n401) );
  INV_X1 U4 ( .A(n407), .ZN(n400) );
  AOI22_X1 U5 ( .A1(n2059), .A2(n408), .B1(n2076), .B2(n409), .ZN(n399) );
  INV_X1 U6 ( .A(n413), .ZN(n398) );
  NAND2_X1 U7 ( .A1(n415), .A2(n417), .ZN(N117) );
  NAND2_X1 U8 ( .A1(n430), .A2(n431), .ZN(N116) );
  AOI21_X1 U9 ( .B1(n2130), .B2(n387), .A(n388), .ZN(n385) );
  NOR2_X1 U10 ( .A1(n1022), .A2(n2144), .ZN(n388) );
  AOI21_X1 U11 ( .B1(n132), .B2(n390), .A(n391), .ZN(n384) );
  NOR2_X1 U12 ( .A1(n1150), .A2(n2099), .ZN(n391) );
  AOI21_X1 U13 ( .B1(n2075), .B2(n393), .A(n394), .ZN(n383) );
  NOR2_X1 U14 ( .A1(n830), .A2(n95), .ZN(n394) );
  AOI21_X1 U15 ( .B1(n2044), .B2(n396), .A(n397), .ZN(n382) );
  NOR2_X1 U16 ( .A1(n894), .A2(n102), .ZN(n397) );
  CLKBUF_X1 U17 ( .A(n130), .Z(n2153) );
  BUF_X2 U18 ( .A(n130), .Z(n2152) );
  INV_X2 U19 ( .A(n2149), .ZN(n2150) );
  INV_X2 U20 ( .A(n2149), .ZN(n2151) );
  BUF_X2 U21 ( .A(n1), .Z(n2192) );
  BUF_X2 U22 ( .A(n2192), .Z(n2194) );
  AND2_X1 U23 ( .A1(n2062), .A2(n2329), .ZN(n1) );
  BUF_X1 U24 ( .A(n121), .Z(n2161) );
  BUF_X2 U25 ( .A(n121), .Z(n2160) );
  INV_X2 U26 ( .A(n109), .ZN(n110) );
  BUF_X2 U27 ( .A(n110), .Z(n2017) );
  BUF_X2 U28 ( .A(n110), .Z(n2016) );
  BUF_X1 U29 ( .A(n109), .Z(n2171) );
  BUF_X2 U30 ( .A(n109), .Z(n2170) );
  CLKBUF_X1 U31 ( .A(n118), .Z(n2162) );
  BUF_X2 U32 ( .A(n118), .Z(n2163) );
  BUF_X1 U33 ( .A(n106), .Z(n2174) );
  BUF_X1 U34 ( .A(n106), .Z(n2172) );
  BUF_X1 U35 ( .A(n106), .Z(n2173) );
  CLKBUF_X3 U36 ( .A(n2), .Z(n2202) );
  CLKBUF_X3 U37 ( .A(n2), .Z(n2201) );
  AND2_X1 U38 ( .A1(n2070), .A2(n2329), .ZN(n2) );
  INV_X2 U39 ( .A(n98), .ZN(n97) );
  BUF_X2 U40 ( .A(n97), .Z(n2025) );
  CLKBUF_X3 U41 ( .A(n98), .Z(n2184) );
  CLKBUF_X3 U42 ( .A(n98), .Z(n2183) );
  BUF_X1 U43 ( .A(n98), .Z(n2182) );
  INV_X2 U44 ( .A(n101), .ZN(n100) );
  BUF_X2 U45 ( .A(n100), .Z(n2024) );
  CLKBUF_X3 U46 ( .A(n101), .Z(n2180) );
  CLKBUF_X3 U47 ( .A(n101), .Z(n2181) );
  BUF_X1 U48 ( .A(n101), .Z(n2179) );
  INV_X2 U49 ( .A(n94), .ZN(n93) );
  BUF_X2 U50 ( .A(n93), .Z(n2026) );
  CLKBUF_X3 U51 ( .A(n94), .Z(n2186) );
  CLKBUF_X3 U52 ( .A(n94), .Z(n2187) );
  BUF_X1 U53 ( .A(n94), .Z(n2185) );
  INV_X2 U54 ( .A(n116), .ZN(n115) );
  BUF_X2 U55 ( .A(n115), .Z(n2014) );
  CLKBUF_X3 U56 ( .A(n116), .Z(n2166) );
  CLKBUF_X3 U57 ( .A(n116), .Z(n2165) );
  BUF_X1 U58 ( .A(n116), .Z(n2164) );
  INV_X2 U59 ( .A(n113), .ZN(n112) );
  BUF_X2 U60 ( .A(n112), .Z(n2015) );
  CLKBUF_X3 U61 ( .A(n113), .Z(n2168) );
  CLKBUF_X3 U62 ( .A(n113), .Z(n2169) );
  BUF_X1 U63 ( .A(n113), .Z(n2167) );
  CLKBUF_X3 U64 ( .A(n128), .Z(n2154) );
  NOR2_X1 U67 ( .A1(CURR_PC[2]), .A2(CURR_PC[3]), .ZN(n697) );
  NOR2_X1 U68 ( .A1(n712), .A2(CURR_PC[2]), .ZN(n694) );
  NOR2_X1 U69 ( .A1(n698), .A2(CURR_PC[5]), .ZN(n693) );
  NOR2_X1 U70 ( .A1(n713), .A2(CURR_PC[3]), .ZN(n696) );
  NOR2_X1 U71 ( .A1(CURR_PC[4]), .A2(CURR_PC[5]), .ZN(n702) );
  BUF_X1 U72 ( .A(n1), .Z(n2191) );
  BUF_X1 U75 ( .A(n103), .Z(n2021) );
  BUF_X1 U76 ( .A(n124), .Z(n2005) );
  BUF_X1 U77 ( .A(n127), .Z(n2003) );
  BUF_X1 U78 ( .A(n2191), .Z(n2195) );
  BUF_X1 U79 ( .A(n2191), .Z(n2193) );
  CLKBUF_X1 U80 ( .A(n104), .Z(n2177) );
  CLKBUF_X1 U81 ( .A(n125), .Z(n2158) );
  INV_X1 U82 ( .A(n2203), .ZN(n2199) );
  INV_X1 U83 ( .A(n2203), .ZN(n2198) );
  BUF_X1 U84 ( .A(n2148), .Z(n1998) );
  CLKBUF_X1 U85 ( .A(n2149), .Z(n1999) );
  CLKBUF_X1 U86 ( .A(n2149), .Z(n1997) );
  INV_X1 U87 ( .A(n2197), .ZN(n2189) );
  INV_X1 U88 ( .A(n2197), .ZN(n2188) );
  BUF_X1 U89 ( .A(n127), .Z(n2004) );
  BUF_X1 U90 ( .A(n103), .Z(n2022) );
  BUF_X1 U91 ( .A(n124), .Z(n2006) );
  BUF_X1 U92 ( .A(n107), .Z(n2019) );
  BUF_X1 U93 ( .A(n119), .Z(n2012) );
  BUF_X1 U94 ( .A(n122), .Z(n2009) );
  CLKBUF_X1 U95 ( .A(n107), .Z(n2018) );
  CLKBUF_X1 U96 ( .A(n119), .Z(n2011) );
  CLKBUF_X1 U97 ( .A(n122), .Z(n2008) );
  CLKBUF_X1 U98 ( .A(n122), .Z(n2010) );
  CLKBUF_X1 U99 ( .A(n107), .Z(n2020) );
  CLKBUF_X1 U100 ( .A(n119), .Z(n2013) );
  CLKBUF_X1 U101 ( .A(n103), .Z(n2023) );
  CLKBUF_X1 U102 ( .A(n124), .Z(n2007) );
  BUF_X1 U103 ( .A(n2), .Z(n2203) );
  BUF_X1 U104 ( .A(n131), .Z(n2001) );
  CLKBUF_X1 U105 ( .A(n131), .Z(n2000) );
  CLKBUF_X1 U106 ( .A(n131), .Z(n2002) );
  BUF_X1 U107 ( .A(n2191), .Z(n2196) );
  BUF_X1 U108 ( .A(n1), .Z(n2197) );
  INV_X1 U109 ( .A(n2178), .ZN(n103) );
  INV_X1 U110 ( .A(n2159), .ZN(n124) );
  INV_X1 U111 ( .A(n2155), .ZN(n127) );
  INV_X1 U112 ( .A(n106), .ZN(n107) );
  INV_X1 U113 ( .A(n118), .ZN(n119) );
  INV_X1 U114 ( .A(n121), .ZN(n122) );
  BUF_X2 U115 ( .A(n128), .Z(n2155) );
  CLKBUF_X1 U116 ( .A(n104), .Z(n2176) );
  CLKBUF_X1 U117 ( .A(n125), .Z(n2157) );
  CLKBUF_X1 U118 ( .A(n104), .Z(n2175) );
  CLKBUF_X1 U119 ( .A(n125), .Z(n2156) );
  BUF_X1 U120 ( .A(n104), .Z(n2178) );
  BUF_X1 U121 ( .A(n125), .Z(n2159) );
  INV_X1 U122 ( .A(n133), .ZN(n2148) );
  INV_X1 U123 ( .A(n133), .ZN(n2149) );
  INV_X1 U124 ( .A(n130), .ZN(n131) );
  NOR2_X1 U127 ( .A1(n2110), .A2(n2366), .ZN(n128) );
  NOR2_X1 U128 ( .A1(n2139), .A2(n2366), .ZN(n113) );
  NOR2_X1 U129 ( .A1(n2053), .A2(n2366), .ZN(n104) );
  NOR2_X1 U130 ( .A1(n2103), .A2(n2366), .ZN(n125) );
  NAND2_X1 U131 ( .A1(n2048), .A2(n2329), .ZN(n106) );
  NAND2_X1 U132 ( .A1(n2125), .A2(n2329), .ZN(n118) );
  NAND2_X1 U133 ( .A1(n2035), .A2(n2329), .ZN(n109) );
  NAND2_X1 U134 ( .A1(n2117), .A2(n2329), .ZN(n121) );
  NAND2_X1 U137 ( .A1(n2088), .A2(n2329), .ZN(n133) );
  BUF_X1 U139 ( .A(n2063), .Z(n2068) );
  BUF_X1 U140 ( .A(n2064), .Z(n2071) );
  BUF_X1 U141 ( .A(n2064), .Z(n2069) );
  BUF_X1 U142 ( .A(n2064), .Z(n2072) );
  BUF_X1 U143 ( .A(n2063), .Z(n2066) );
  BUF_X1 U144 ( .A(n2063), .Z(n2067) );
  BUF_X1 U145 ( .A(n2063), .Z(n2065) );
  BUF_X1 U146 ( .A(n136), .Z(n2073) );
  BUF_X1 U147 ( .A(n136), .Z(n2074) );
  BUF_X1 U148 ( .A(n2064), .Z(n2070) );
  BUF_X1 U149 ( .A(n136), .Z(n2075) );
  BUF_X1 U150 ( .A(n136), .Z(n2076) );
  INV_X1 U151 ( .A(n12), .ZN(n11) );
  INV_X1 U152 ( .A(n14), .ZN(n13) );
  BUF_X1 U153 ( .A(n2204), .Z(n2214) );
  BUF_X1 U154 ( .A(n2204), .Z(n2215) );
  NOR2_X1 U155 ( .A1(n2146), .A2(n2366), .ZN(n116) );
  NOR2_X1 U156 ( .A1(n2077), .A2(n2366), .ZN(n94) );
  NOR2_X1 U157 ( .A1(n2049), .A2(n2366), .ZN(n101) );
  NOR2_X1 U158 ( .A1(n2079), .A2(n2366), .ZN(n98) );
  NAND2_X1 U159 ( .A1(n2095), .A2(n2329), .ZN(n130) );
  BUF_X1 U161 ( .A(n105), .Z(n2054) );
  BUF_X1 U162 ( .A(n105), .Z(n2052) );
  BUF_X1 U163 ( .A(n105), .Z(n2051) );
  BUF_X1 U164 ( .A(n105), .Z(n2053) );
  BUF_X1 U165 ( .A(n2097), .Z(n2098) );
  BUF_X1 U166 ( .A(n126), .Z(n2101) );
  BUF_X1 U167 ( .A(n2097), .Z(n2099) );
  BUF_X1 U168 ( .A(n2097), .Z(n2100) );
  BUF_X1 U169 ( .A(n105), .Z(n2055) );
  BUF_X1 U170 ( .A(n2132), .Z(n2135) );
  BUF_X1 U171 ( .A(n2132), .Z(n2134) );
  BUF_X1 U172 ( .A(n2132), .Z(n2136) );
  BUF_X1 U173 ( .A(n2132), .Z(n2137) );
  BUF_X1 U174 ( .A(n2133), .Z(n2141) );
  BUF_X1 U175 ( .A(n2133), .Z(n2140) );
  BUF_X1 U176 ( .A(n2133), .Z(n2138) );
  BUF_X1 U177 ( .A(n114), .Z(n2142) );
  BUF_X1 U178 ( .A(n114), .Z(n2143) );
  BUF_X1 U179 ( .A(n2104), .Z(n2105) );
  BUF_X1 U180 ( .A(n129), .Z(n2108) );
  BUF_X1 U181 ( .A(n2104), .Z(n2106) );
  BUF_X1 U182 ( .A(n2104), .Z(n2107) );
  BUF_X1 U183 ( .A(n2133), .Z(n2139) );
  AND2_X1 U184 ( .A1(n706), .A2(n695), .ZN(n2063) );
  AND2_X1 U185 ( .A1(n706), .A2(n695), .ZN(n2064) );
  BUF_X1 U186 ( .A(n123), .Z(n2115) );
  BUF_X1 U187 ( .A(n2111), .Z(n2113) );
  BUF_X1 U188 ( .A(n2111), .Z(n2114) );
  BUF_X1 U189 ( .A(n2111), .Z(n2112) );
  BUF_X1 U190 ( .A(n91), .Z(n2060) );
  BUF_X1 U191 ( .A(n2056), .Z(n2058) );
  BUF_X1 U192 ( .A(n2056), .Z(n2059) );
  BUF_X1 U193 ( .A(n2056), .Z(n2057) );
  BUF_X1 U194 ( .A(n2081), .Z(n2084) );
  BUF_X1 U195 ( .A(n2081), .Z(n2085) );
  BUF_X1 U196 ( .A(n2081), .Z(n2086) );
  BUF_X1 U197 ( .A(n2082), .Z(n2090) );
  BUF_X1 U198 ( .A(n2082), .Z(n2089) );
  BUF_X1 U199 ( .A(n2082), .Z(n2087) );
  BUF_X1 U200 ( .A(n2081), .Z(n2083) );
  BUF_X1 U201 ( .A(n2028), .Z(n2031) );
  BUF_X1 U202 ( .A(n2028), .Z(n2032) );
  BUF_X1 U203 ( .A(n2028), .Z(n2033) );
  BUF_X1 U204 ( .A(n2029), .Z(n2036) );
  BUF_X1 U205 ( .A(n2029), .Z(n2034) );
  BUF_X1 U206 ( .A(n2029), .Z(n2037) );
  BUF_X1 U207 ( .A(n2028), .Z(n2030) );
  BUF_X1 U208 ( .A(n135), .Z(n2091) );
  BUF_X1 U209 ( .A(n135), .Z(n2092) );
  AND2_X1 U210 ( .A1(n706), .A2(n695), .ZN(n136) );
  BUF_X1 U211 ( .A(n111), .Z(n2038) );
  BUF_X1 U212 ( .A(n111), .Z(n2039) );
  BUF_X1 U213 ( .A(n2042), .Z(n2045) );
  BUF_X1 U214 ( .A(n108), .Z(n2046) );
  BUF_X1 U215 ( .A(n2042), .Z(n2044) );
  BUF_X1 U216 ( .A(n2042), .Z(n2043) );
  BUF_X1 U217 ( .A(n2082), .Z(n2088) );
  BUF_X1 U218 ( .A(n2029), .Z(n2035) );
  BUF_X1 U219 ( .A(n2118), .Z(n2123) );
  BUF_X1 U220 ( .A(n2119), .Z(n2126) );
  BUF_X1 U221 ( .A(n2119), .Z(n2124) );
  BUF_X1 U222 ( .A(n2119), .Z(n2127) );
  BUF_X1 U223 ( .A(n2118), .Z(n2121) );
  BUF_X1 U224 ( .A(n2118), .Z(n2122) );
  BUF_X1 U225 ( .A(n2118), .Z(n2120) );
  BUF_X1 U226 ( .A(n120), .Z(n2128) );
  BUF_X1 U227 ( .A(n120), .Z(n2129) );
  BUF_X1 U228 ( .A(n2119), .Z(n2125) );
  BUF_X1 U229 ( .A(n126), .Z(n2102) );
  BUF_X1 U230 ( .A(n126), .Z(n2103) );
  BUF_X1 U231 ( .A(n129), .Z(n2109) );
  BUF_X1 U232 ( .A(n129), .Z(n2110) );
  BUF_X1 U233 ( .A(n123), .Z(n2116) );
  BUF_X1 U234 ( .A(n91), .Z(n2061) );
  BUF_X1 U235 ( .A(n123), .Z(n2117) );
  BUF_X1 U236 ( .A(n91), .Z(n2062) );
  BUF_X1 U237 ( .A(n108), .Z(n2047) );
  BUF_X1 U238 ( .A(n108), .Z(n2048) );
  AND2_X1 U239 ( .A1(n2325), .A2(n2324), .ZN(n1964) );
  BUF_X1 U240 ( .A(n135), .Z(n2093) );
  BUF_X1 U241 ( .A(n111), .Z(n2040) );
  BUF_X1 U242 ( .A(n120), .Z(n2130) );
  BUF_X1 U244 ( .A(n114), .Z(n2144) );
  BUF_X1 U245 ( .A(n114), .Z(n2145) );
  BUF_X1 U246 ( .A(n135), .Z(n2094) );
  BUF_X1 U247 ( .A(n111), .Z(n2041) );
  BUF_X1 U248 ( .A(n120), .Z(n2131) );
  NAND2_X1 U249 ( .A1(n45), .A2(n46), .ZN(n12) );
  NAND2_X1 U250 ( .A1(n45), .A2(n47), .ZN(n14) );
  INV_X1 U251 ( .A(n10), .ZN(n8) );
  INV_X1 U252 ( .A(n16), .ZN(n15) );
  INV_X1 U253 ( .A(n18), .ZN(n17) );
  INV_X1 U254 ( .A(n20), .ZN(n19) );
  INV_X1 U255 ( .A(n22), .ZN(n21) );
  INV_X1 U256 ( .A(n24), .ZN(n23) );
  INV_X1 U257 ( .A(n26), .ZN(n25) );
  INV_X1 U258 ( .A(n28), .ZN(n27) );
  INV_X1 U259 ( .A(n30), .ZN(n29) );
  INV_X1 U260 ( .A(n32), .ZN(n31) );
  INV_X1 U261 ( .A(n34), .ZN(n33) );
  INV_X1 U262 ( .A(n36), .ZN(n35) );
  INV_X1 U263 ( .A(n38), .ZN(n37) );
  INV_X1 U264 ( .A(n40), .ZN(n39) );
  BUF_X1 U265 ( .A(RST), .Z(n2204) );
  NOR2_X1 U266 ( .A1(n712), .A2(n713), .ZN(n695) );
  NOR2_X1 U267 ( .A1(n707), .A2(n698), .ZN(n706) );
  MUX2_X1 U268 ( .A(n2218), .B(n2220), .S(n2219), .Z(n2328) );
  MUX2_X1 U269 ( .A(N850), .B(n2220), .S(n2219), .Z(n2327) );
  NAND2_X1 U270 ( .A1(n711), .A2(n695), .ZN(n2049) );
  NAND2_X1 U271 ( .A1(n696), .A2(n706), .ZN(n2077) );
  NAND2_X1 U272 ( .A1(n693), .A2(n694), .ZN(n2146) );
  NAND2_X1 U273 ( .A1(n697), .A2(n706), .ZN(n2079) );
  NAND2_X1 U274 ( .A1(n711), .A2(n695), .ZN(n102) );
  NAND2_X1 U275 ( .A1(n711), .A2(n695), .ZN(n2050) );
  NAND2_X1 U276 ( .A1(n696), .A2(n706), .ZN(n95) );
  NAND2_X1 U277 ( .A1(n696), .A2(n706), .ZN(n2078) );
  NAND2_X1 U278 ( .A1(n693), .A2(n694), .ZN(n117) );
  NAND2_X1 U279 ( .A1(n693), .A2(n694), .ZN(n2147) );
  NAND2_X1 U280 ( .A1(n697), .A2(n706), .ZN(n99) );
  NAND2_X1 U281 ( .A1(n697), .A2(n706), .ZN(n2080) );
  AND2_X1 U282 ( .A1(n702), .A2(n696), .ZN(n132) );
  AND2_X1 U283 ( .A1(n702), .A2(n696), .ZN(n2096) );
  NAND2_X1 U284 ( .A1(n711), .A2(n694), .ZN(n105) );
  AND2_X1 U285 ( .A1(n702), .A2(n696), .ZN(n2095) );
  NAND2_X1 U286 ( .A1(n702), .A2(n695), .ZN(n126) );
  NAND2_X1 U287 ( .A1(n702), .A2(n694), .ZN(n129) );
  NAND2_X1 U288 ( .A1(n702), .A2(n695), .ZN(n2097) );
  NAND2_X1 U289 ( .A1(n702), .A2(n694), .ZN(n2104) );
  NAND2_X1 U290 ( .A1(n693), .A2(n695), .ZN(n2132) );
  NAND2_X1 U291 ( .A1(n693), .A2(n695), .ZN(n2133) );
  NAND2_X1 U292 ( .A1(n693), .A2(n695), .ZN(n114) );
  NAND4_X1 U293 ( .A1(n366), .A2(n367), .A3(n368), .A4(n369), .ZN(N120) );
  AOI221_X1 U294 ( .B1(n2057), .B2(n376), .C1(n2074), .C2(n377), .A(n378), 
        .ZN(n367) );
  AOI221_X1 U295 ( .B1(n2112), .B2(n370), .C1(n2129), .C2(n371), .A(n372), 
        .ZN(n369) );
  AOI221_X1 U296 ( .B1(n2039), .B2(n379), .C1(n2043), .C2(n380), .A(n381), 
        .ZN(n366) );
  NAND4_X1 U297 ( .A1(n334), .A2(n335), .A3(n336), .A4(n337), .ZN(N90) );
  AOI221_X1 U298 ( .B1(n2060), .B2(n344), .C1(n2072), .C2(n345), .A(n346), 
        .ZN(n335) );
  AOI221_X1 U299 ( .B1(n2115), .B2(n338), .C1(n2127), .C2(n339), .A(n340), 
        .ZN(n337) );
  AOI221_X1 U300 ( .B1(n2037), .B2(n347), .C1(n2046), .C2(n348), .A(n349), 
        .ZN(n334) );
  NOR3_X1 U301 ( .A1(INST_29), .A2(INST_31), .A3(INST_30), .ZN(n715) );
  NAND4_X1 U302 ( .A1(n686), .A2(n687), .A3(n688), .A4(n689), .ZN(N100) );
  AOI221_X1 U303 ( .B1(n2117), .B2(n690), .C1(n2122), .C2(n691), .A(n692), 
        .ZN(n689) );
  AOI221_X1 U304 ( .B1(n2062), .B2(n703), .C1(n2067), .C2(n704), .A(n705), 
        .ZN(n687) );
  AOI221_X1 U305 ( .B1(n2032), .B2(n708), .C1(n2048), .C2(n709), .A(n710), 
        .ZN(n686) );
  NAND4_X1 U306 ( .A1(n670), .A2(n671), .A3(n672), .A4(n673), .ZN(N101) );
  AOI221_X1 U307 ( .B1(n2061), .B2(n680), .C1(n2066), .C2(n681), .A(n682), 
        .ZN(n671) );
  AOI221_X1 U308 ( .B1(n2116), .B2(n674), .C1(n2121), .C2(n675), .A(n676), 
        .ZN(n673) );
  AOI221_X1 U309 ( .B1(n2031), .B2(n683), .C1(n2047), .C2(n684), .A(n685), 
        .ZN(n670) );
  NAND4_X1 U310 ( .A1(n654), .A2(n655), .A3(n656), .A4(n657), .ZN(N102) );
  AOI221_X1 U311 ( .B1(n2060), .B2(n664), .C1(n2065), .C2(n665), .A(n666), 
        .ZN(n655) );
  AOI221_X1 U312 ( .B1(n2115), .B2(n658), .C1(n2120), .C2(n659), .A(n660), 
        .ZN(n657) );
  AOI221_X1 U313 ( .B1(n2030), .B2(n667), .C1(n2046), .C2(n668), .A(n669), 
        .ZN(n654) );
  NAND4_X1 U314 ( .A1(n238), .A2(n239), .A3(n240), .A4(n241), .ZN(N96) );
  AOI221_X1 U315 ( .B1(n2058), .B2(n248), .C1(n2069), .C2(n249), .A(n250), 
        .ZN(n239) );
  AOI221_X1 U316 ( .B1(n2113), .B2(n242), .C1(n2124), .C2(n243), .A(n244), 
        .ZN(n241) );
  AOI221_X1 U317 ( .B1(n2034), .B2(n251), .C1(n2044), .C2(n252), .A(n253), 
        .ZN(n238) );
  NAND4_X1 U318 ( .A1(n222), .A2(n223), .A3(n224), .A4(n225), .ZN(N97) );
  AOI221_X1 U319 ( .B1(n2057), .B2(n232), .C1(n2068), .C2(n233), .A(n234), 
        .ZN(n223) );
  AOI221_X1 U320 ( .B1(n2112), .B2(n226), .C1(n2123), .C2(n227), .A(n228), 
        .ZN(n225) );
  AOI221_X1 U321 ( .B1(n2033), .B2(n235), .C1(n2043), .C2(n236), .A(n237), 
        .ZN(n222) );
  NAND4_X1 U322 ( .A1(n206), .A2(n207), .A3(n208), .A4(n209), .ZN(N98) );
  AOI221_X1 U323 ( .B1(n2114), .B2(n210), .C1(n2122), .C2(n211), .A(n212), 
        .ZN(n209) );
  AOI221_X1 U324 ( .B1(n2059), .B2(n216), .C1(n2067), .C2(n217), .A(n218), 
        .ZN(n207) );
  AOI221_X1 U325 ( .B1(n2032), .B2(n219), .C1(n2045), .C2(n220), .A(n221), 
        .ZN(n206) );
  NAND4_X1 U326 ( .A1(n302), .A2(n303), .A3(n304), .A4(n305), .ZN(N92) );
  AOI221_X1 U327 ( .B1(n2117), .B2(n306), .C1(n2128), .C2(n307), .A(n308), 
        .ZN(n305) );
  AOI221_X1 U328 ( .B1(n2062), .B2(n312), .C1(n2073), .C2(n313), .A(n314), 
        .ZN(n303) );
  AOI221_X1 U329 ( .B1(n2038), .B2(n315), .C1(n2048), .C2(n316), .A(n317), 
        .ZN(n302) );
  NAND4_X1 U330 ( .A1(n286), .A2(n287), .A3(n288), .A4(n289), .ZN(N93) );
  AOI221_X1 U331 ( .B1(n2061), .B2(n296), .C1(n2072), .C2(n297), .A(n298), 
        .ZN(n287) );
  AOI221_X1 U332 ( .B1(n2116), .B2(n290), .C1(n2127), .C2(n291), .A(n292), 
        .ZN(n289) );
  AOI221_X1 U333 ( .B1(n2037), .B2(n299), .C1(n2047), .C2(n300), .A(n301), 
        .ZN(n286) );
  NAND4_X1 U334 ( .A1(n270), .A2(n271), .A3(n272), .A4(n273), .ZN(N94) );
  AOI221_X1 U335 ( .B1(n2060), .B2(n280), .C1(n2071), .C2(n281), .A(n282), 
        .ZN(n271) );
  AOI221_X1 U336 ( .B1(n2115), .B2(n274), .C1(n2126), .C2(n275), .A(n276), 
        .ZN(n273) );
  AOI221_X1 U337 ( .B1(n2036), .B2(n283), .C1(n2046), .C2(n284), .A(n285), 
        .ZN(n270) );
  NAND4_X1 U338 ( .A1(n638), .A2(n639), .A3(n640), .A4(n641), .ZN(N103) );
  AOI221_X1 U339 ( .B1(n2116), .B2(n642), .C1(n2131), .C2(n643), .A(n644), 
        .ZN(n641) );
  AOI221_X1 U340 ( .B1(n2061), .B2(n648), .C1(n2076), .C2(n649), .A(n650), 
        .ZN(n639) );
  AOI221_X1 U341 ( .B1(n2041), .B2(n651), .C1(n2047), .C2(n652), .A(n653), 
        .ZN(n638) );
  NAND4_X1 U342 ( .A1(n606), .A2(n607), .A3(n608), .A4(n609), .ZN(N105) );
  AOI221_X1 U343 ( .B1(n2059), .B2(n616), .C1(n2074), .C2(n617), .A(n618), 
        .ZN(n607) );
  AOI221_X1 U344 ( .B1(n2114), .B2(n610), .C1(n2129), .C2(n611), .A(n612), 
        .ZN(n609) );
  AOI221_X1 U345 ( .B1(n2039), .B2(n619), .C1(n2045), .C2(n620), .A(n621), 
        .ZN(n606) );
  NAND4_X1 U346 ( .A1(n590), .A2(n591), .A3(n592), .A4(n593), .ZN(N106) );
  AOI221_X1 U347 ( .B1(n2114), .B2(n594), .C1(n2128), .C2(n595), .A(n596), 
        .ZN(n593) );
  AOI221_X1 U348 ( .B1(n2059), .B2(n600), .C1(n2073), .C2(n601), .A(n602), 
        .ZN(n591) );
  AOI221_X1 U349 ( .B1(n2038), .B2(n603), .C1(n2045), .C2(n604), .A(n605), 
        .ZN(n590) );
  NAND4_X1 U350 ( .A1(n494), .A2(n495), .A3(n496), .A4(n497), .ZN(N112) );
  AOI221_X1 U351 ( .B1(n2117), .B2(n498), .C1(n2125), .C2(n499), .A(n500), 
        .ZN(n497) );
  AOI221_X1 U352 ( .B1(n2062), .B2(n504), .C1(n2070), .C2(n505), .A(n506), 
        .ZN(n495) );
  AOI221_X1 U353 ( .B1(n2035), .B2(n507), .C1(n2048), .C2(n508), .A(n509), 
        .ZN(n494) );
  NAND4_X1 U354 ( .A1(n478), .A2(n479), .A3(n480), .A4(n481), .ZN(N113) );
  AOI221_X1 U355 ( .B1(n2061), .B2(n488), .C1(n2069), .C2(n489), .A(n490), 
        .ZN(n479) );
  AOI221_X1 U356 ( .B1(n2116), .B2(n482), .C1(n2124), .C2(n483), .A(n484), 
        .ZN(n481) );
  AOI221_X1 U357 ( .B1(n2034), .B2(n491), .C1(n2047), .C2(n492), .A(n493), 
        .ZN(n478) );
  NAND4_X1 U358 ( .A1(n462), .A2(n463), .A3(n464), .A4(n465), .ZN(N114) );
  AOI221_X1 U359 ( .B1(n2060), .B2(n472), .C1(n2068), .C2(n473), .A(n474), 
        .ZN(n463) );
  AOI221_X1 U360 ( .B1(n2115), .B2(n466), .C1(n2123), .C2(n467), .A(n468), 
        .ZN(n465) );
  AOI221_X1 U361 ( .B1(n2033), .B2(n475), .C1(n2046), .C2(n476), .A(n477), 
        .ZN(n462) );
  NAND4_X1 U362 ( .A1(n558), .A2(n559), .A3(n560), .A4(n561), .ZN(N108) );
  AOI221_X1 U363 ( .B1(n2057), .B2(n568), .C1(n2071), .C2(n569), .A(n570), 
        .ZN(n559) );
  AOI221_X1 U364 ( .B1(n2112), .B2(n562), .C1(n2126), .C2(n563), .A(n564), 
        .ZN(n561) );
  AOI221_X1 U365 ( .B1(n2036), .B2(n571), .C1(n2043), .C2(n572), .A(n573), 
        .ZN(n558) );
  NAND4_X1 U366 ( .A1(n542), .A2(n543), .A3(n544), .A4(n545), .ZN(N109) );
  AOI221_X1 U367 ( .B1(n2115), .B2(n546), .C1(n2124), .C2(n547), .A(n548), 
        .ZN(n545) );
  AOI221_X1 U368 ( .B1(n2060), .B2(n552), .C1(n2069), .C2(n553), .A(n554), 
        .ZN(n543) );
  AOI221_X1 U369 ( .B1(n2034), .B2(n555), .C1(n2046), .C2(n556), .A(n557), 
        .ZN(n542) );
  NAND4_X1 U370 ( .A1(n526), .A2(n527), .A3(n528), .A4(n529), .ZN(N110) );
  AOI221_X1 U371 ( .B1(n2058), .B2(n536), .C1(n2074), .C2(n537), .A(n538), 
        .ZN(n527) );
  AOI221_X1 U372 ( .B1(n2113), .B2(n530), .C1(n2129), .C2(n531), .A(n532), 
        .ZN(n529) );
  AOI221_X1 U373 ( .B1(n2039), .B2(n539), .C1(n2044), .C2(n540), .A(n541), 
        .ZN(n526) );
  AND2_X1 U374 ( .A1(n693), .A2(n697), .ZN(n123) );
  AND2_X1 U375 ( .A1(n693), .A2(n697), .ZN(n2111) );
  AND2_X1 U376 ( .A1(n694), .A2(n706), .ZN(n91) );
  AND2_X1 U377 ( .A1(n694), .A2(n706), .ZN(n2056) );
  AND2_X1 U378 ( .A1(n711), .A2(n696), .ZN(n2042) );
  AND2_X1 U379 ( .A1(n711), .A2(n696), .ZN(n108) );
  AND2_X1 U380 ( .A1(n693), .A2(n696), .ZN(n2118) );
  AND2_X1 U381 ( .A1(n693), .A2(n696), .ZN(n2119) );
  AND2_X1 U382 ( .A1(n702), .A2(n697), .ZN(n2081) );
  AND2_X1 U383 ( .A1(n702), .A2(n697), .ZN(n2082) );
  AND2_X1 U384 ( .A1(n693), .A2(n696), .ZN(n120) );
  AND2_X1 U385 ( .A1(n711), .A2(n697), .ZN(n2028) );
  AND2_X1 U386 ( .A1(n711), .A2(n697), .ZN(n2029) );
  AND2_X1 U387 ( .A1(n702), .A2(n697), .ZN(n135) );
  AND2_X1 U388 ( .A1(n711), .A2(n697), .ZN(n111) );
  NAND4_X1 U389 ( .A1(n350), .A2(n351), .A3(n352), .A4(n353), .ZN(N121) );
  AOI221_X1 U390 ( .B1(n2113), .B2(n354), .C1(n2123), .C2(n355), .A(n356), 
        .ZN(n353) );
  AOI221_X1 U391 ( .B1(n2058), .B2(n360), .C1(n2068), .C2(n361), .A(n362), 
        .ZN(n351) );
  NOR2_X1 U392 ( .A1(\PC_HISTORY[1][2] ), .A2(\PC_HISTORY[1][3] ), .ZN(n45) );
  AOI221_X1 U393 ( .B1(n2112), .B2(\PRED_TABLE[4][1] ), .C1(n2120), .C2(
        \PRED_TABLE[5][1] ), .A(n180), .ZN(n177) );
  AOI221_X1 U394 ( .B1(n2057), .B2(\PRED_TABLE[14][1] ), .C1(n2065), .C2(
        \PRED_TABLE[15][1] ), .A(n186), .ZN(n175) );
  AOI221_X1 U395 ( .B1(n2083), .B2(\PRED_TABLE[0][1] ), .C1(n2096), .C2(
        \PRED_TABLE[1][1] ), .A(n183), .ZN(n176) );
  AND2_X1 U396 ( .A1(n57), .A2(\PC_HISTORY[1][0] ), .ZN(n47) );
  AND2_X1 U397 ( .A1(n51), .A2(\PC_HISTORY[1][0] ), .ZN(n46) );
  NAND2_X1 U398 ( .A1(n50), .A2(n47), .ZN(n10) );
  NAND2_X1 U399 ( .A1(n48), .A2(n46), .ZN(n16) );
  NAND2_X1 U400 ( .A1(n48), .A2(n47), .ZN(n18) );
  NAND2_X1 U401 ( .A1(n49), .A2(n46), .ZN(n20) );
  NAND2_X1 U402 ( .A1(n49), .A2(n47), .ZN(n22) );
  NAND2_X1 U403 ( .A1(n46), .A2(n50), .ZN(n24) );
  NAND2_X1 U404 ( .A1(n53), .A2(n50), .ZN(n26) );
  NAND2_X1 U405 ( .A1(n54), .A2(n50), .ZN(n28) );
  NAND2_X1 U406 ( .A1(n53), .A2(n49), .ZN(n30) );
  NAND2_X1 U407 ( .A1(n54), .A2(n49), .ZN(n32) );
  NAND2_X1 U408 ( .A1(n53), .A2(n48), .ZN(n34) );
  NAND2_X1 U409 ( .A1(n54), .A2(n48), .ZN(n36) );
  NAND2_X1 U410 ( .A1(n53), .A2(n45), .ZN(n38) );
  NAND2_X1 U411 ( .A1(n54), .A2(n45), .ZN(n40) );
  NOR2_X1 U412 ( .A1(n707), .A2(CURR_PC[4]), .ZN(n711) );
  AOI221_X1 U413 ( .B1(n2086), .B2(n357), .C1(n2095), .C2(n358), .A(n359), 
        .ZN(n352) );
  OAI22_X1 U414 ( .A1(n1151), .A2(n2099), .B1(n1183), .B2(n2106), .ZN(n359) );
  AOI221_X1 U415 ( .B1(n2084), .B2(n197), .C1(n132), .C2(n198), .A(n199), .ZN(
        n192) );
  OAI22_X1 U416 ( .A1(n1140), .A2(n2099), .B1(n1172), .B2(n2106), .ZN(n199) );
  AOI221_X1 U417 ( .B1(n2085), .B2(n699), .C1(n2095), .C2(n700), .A(n701), 
        .ZN(n688) );
  OAI22_X1 U418 ( .A1(n1162), .A2(n2103), .B1(n1194), .B2(n2110), .ZN(n701) );
  AOI221_X1 U419 ( .B1(n2084), .B2(n677), .C1(n132), .C2(n678), .A(n679), .ZN(
        n672) );
  OAI22_X1 U420 ( .A1(n1141), .A2(n2102), .B1(n1173), .B2(n2109), .ZN(n679) );
  AOI221_X1 U421 ( .B1(n2083), .B2(n661), .C1(n2096), .C2(n662), .A(n663), 
        .ZN(n656) );
  OAI22_X1 U422 ( .A1(n1161), .A2(n2101), .B1(n1193), .B2(n2108), .ZN(n663) );
  AOI221_X1 U423 ( .B1(n2088), .B2(n261), .C1(n2095), .C2(n262), .A(n263), 
        .ZN(n256) );
  OAI22_X1 U424 ( .A1(n1138), .A2(n2098), .B1(n1170), .B2(n2105), .ZN(n263) );
  AOI221_X1 U425 ( .B1(n2087), .B2(n245), .C1(n132), .C2(n246), .A(n247), .ZN(
        n240) );
  OAI22_X1 U426 ( .A1(n1164), .A2(n2099), .B1(n1196), .B2(n2106), .ZN(n247) );
  AOI221_X1 U427 ( .B1(n2086), .B2(n229), .C1(n2096), .C2(n230), .A(n231), 
        .ZN(n224) );
  OAI22_X1 U428 ( .A1(n1139), .A2(n2098), .B1(n1171), .B2(n2105), .ZN(n231) );
  AOI221_X1 U429 ( .B1(n2085), .B2(n213), .C1(n2095), .C2(n214), .A(n215), 
        .ZN(n208) );
  OAI22_X1 U430 ( .A1(n1163), .A2(n2100), .B1(n1195), .B2(n2107), .ZN(n215) );
  AOI221_X1 U431 ( .B1(n2089), .B2(n325), .C1(n2096), .C2(n326), .A(n327), 
        .ZN(n320) );
  OAI22_X1 U432 ( .A1(n1136), .A2(n2100), .B1(n1168), .B2(n2107), .ZN(n327) );
  AOI221_X1 U433 ( .B1(n2091), .B2(n309), .C1(n2095), .C2(n310), .A(n311), 
        .ZN(n304) );
  OAI22_X1 U434 ( .A1(n1166), .A2(n2103), .B1(n1198), .B2(n2110), .ZN(n311) );
  AOI221_X1 U435 ( .B1(n2090), .B2(n293), .C1(n132), .C2(n294), .A(n295), .ZN(
        n288) );
  OAI22_X1 U436 ( .A1(n1137), .A2(n2102), .B1(n1169), .B2(n2109), .ZN(n295) );
  AOI221_X1 U437 ( .B1(n2089), .B2(n277), .C1(n2096), .C2(n278), .A(n279), 
        .ZN(n272) );
  OAI22_X1 U438 ( .A1(n1165), .A2(n2101), .B1(n1197), .B2(n2108), .ZN(n279) );
  AOI221_X1 U439 ( .B1(n2093), .B2(n629), .C1(n132), .C2(n630), .A(n631), .ZN(
        n624) );
  OAI22_X1 U440 ( .A1(n1160), .A2(n2101), .B1(n1192), .B2(n2108), .ZN(n631) );
  AOI221_X1 U441 ( .B1(n2094), .B2(n645), .C1(n2095), .C2(n646), .A(n647), 
        .ZN(n640) );
  OAI22_X1 U442 ( .A1(n1142), .A2(n2102), .B1(n1174), .B2(n2109), .ZN(n647) );
  AOI221_X1 U443 ( .B1(n2092), .B2(n613), .C1(n2096), .C2(n614), .A(n615), 
        .ZN(n608) );
  OAI22_X1 U444 ( .A1(n1143), .A2(n2100), .B1(n1175), .B2(n2107), .ZN(n615) );
  AOI221_X1 U445 ( .B1(n2091), .B2(n597), .C1(n2095), .C2(n598), .A(n599), 
        .ZN(n592) );
  OAI22_X1 U446 ( .A1(n1159), .A2(n2100), .B1(n1191), .B2(n2107), .ZN(n599) );
  AOI221_X1 U447 ( .B1(n2091), .B2(n517), .C1(n2096), .C2(n518), .A(n519), 
        .ZN(n512) );
  OAI22_X1 U448 ( .A1(n1146), .A2(n2098), .B1(n1178), .B2(n2105), .ZN(n519) );
  AOI221_X1 U449 ( .B1(n2088), .B2(n501), .C1(n2095), .C2(n502), .A(n503), 
        .ZN(n496) );
  OAI22_X1 U450 ( .A1(n1156), .A2(n2103), .B1(n1188), .B2(n2110), .ZN(n503) );
  AOI221_X1 U451 ( .B1(n2087), .B2(n485), .C1(n132), .C2(n486), .A(n487), .ZN(
        n480) );
  OAI22_X1 U452 ( .A1(n1147), .A2(n2102), .B1(n1179), .B2(n2109), .ZN(n487) );
  AOI221_X1 U453 ( .B1(n2086), .B2(n469), .C1(n2096), .C2(n470), .A(n471), 
        .ZN(n464) );
  OAI22_X1 U454 ( .A1(n1155), .A2(n2101), .B1(n1187), .B2(n2108), .ZN(n471) );
  AOI221_X1 U455 ( .B1(n2090), .B2(n581), .C1(n132), .C2(n582), .A(n583), .ZN(
        n576) );
  OAI22_X1 U456 ( .A1(n1144), .A2(n2099), .B1(n1176), .B2(n2106), .ZN(n583) );
  AOI221_X1 U457 ( .B1(n2089), .B2(n565), .C1(n2096), .C2(n566), .A(n567), 
        .ZN(n560) );
  OAI22_X1 U458 ( .A1(n1158), .A2(n2098), .B1(n1190), .B2(n2105), .ZN(n567) );
  AOI221_X1 U459 ( .B1(n2087), .B2(n549), .C1(n2095), .C2(n550), .A(n551), 
        .ZN(n544) );
  OAI22_X1 U460 ( .A1(n1145), .A2(n2101), .B1(n1177), .B2(n2108), .ZN(n551) );
  AOI221_X1 U461 ( .B1(n2092), .B2(n533), .C1(n132), .C2(n534), .A(n535), .ZN(
        n528) );
  OAI22_X1 U462 ( .A1(n1157), .A2(n2099), .B1(n1189), .B2(n2106), .ZN(n535) );
  AOI221_X1 U463 ( .B1(n2092), .B2(n373), .C1(n2096), .C2(n374), .A(n375), 
        .ZN(n368) );
  OAI22_X1 U464 ( .A1(n1152), .A2(n2098), .B1(n1184), .B2(n2105), .ZN(n375) );
  AOI221_X1 U465 ( .B1(n2090), .B2(n341), .C1(n132), .C2(n342), .A(n343), .ZN(
        n336) );
  OAI22_X1 U466 ( .A1(n1167), .A2(n2101), .B1(n1199), .B2(n2108), .ZN(n343) );
  OAI22_X1 U467 ( .A1(n1153), .A2(n2100), .B1(n1185), .B2(n2107), .ZN(n407) );
  AOI221_X1 U468 ( .B1(n2085), .B2(n453), .C1(n2095), .C2(n454), .A(n455), 
        .ZN(n448) );
  OAI22_X1 U469 ( .A1(n1148), .A2(n2100), .B1(n1180), .B2(n2107), .ZN(n455) );
  AOI221_X1 U470 ( .B1(n2033), .B2(n363), .C1(n2044), .C2(n364), .A(n365), 
        .ZN(n350) );
  OAI22_X1 U471 ( .A1(n895), .A2(n2049), .B1(n927), .B2(n2053), .ZN(n365) );
  AOI221_X1 U472 ( .B1(n2035), .B2(n267), .C1(n2043), .C2(n268), .A(n269), 
        .ZN(n254) );
  OAI22_X1 U473 ( .A1(n882), .A2(n2049), .B1(n914), .B2(n2054), .ZN(n269) );
  OAI22_X1 U474 ( .A1(n897), .A2(n2049), .B1(n929), .B2(n2054), .ZN(n413) );
  AOI221_X1 U475 ( .B1(n2032), .B2(n459), .C1(n2045), .C2(n460), .A(n461), 
        .ZN(n446) );
  OAI22_X1 U476 ( .A1(n892), .A2(n2049), .B1(n924), .B2(n2052), .ZN(n461) );
  AOI221_X1 U477 ( .B1(n2031), .B2(n203), .C1(n2044), .C2(n204), .A(n205), 
        .ZN(n190) );
  OAI22_X1 U478 ( .A1(n884), .A2(n102), .B1(n916), .B2(n2052), .ZN(n205) );
  AOI221_X1 U479 ( .B1(n2036), .B2(n331), .C1(n2045), .C2(n332), .A(n333), 
        .ZN(n318) );
  OAI22_X1 U480 ( .A1(n880), .A2(n2050), .B1(n912), .B2(n2053), .ZN(n333) );
  AOI221_X1 U481 ( .B1(n2040), .B2(n635), .C1(n2046), .C2(n636), .A(n637), 
        .ZN(n622) );
  OAI22_X1 U482 ( .A1(n904), .A2(n102), .B1(n936), .B2(n2054), .ZN(n637) );
  AOI221_X1 U483 ( .B1(n2038), .B2(n523), .C1(n2043), .C2(n524), .A(n525), 
        .ZN(n510) );
  OAI22_X1 U484 ( .A1(n890), .A2(n2050), .B1(n922), .B2(n2054), .ZN(n525) );
  AOI221_X1 U485 ( .B1(n2037), .B2(n587), .C1(n2044), .C2(n588), .A(n589), 
        .ZN(n574) );
  OAI22_X1 U486 ( .A1(n888), .A2(n102), .B1(n920), .B2(n2051), .ZN(n589) );
  AOI221_X1 U487 ( .B1(n2031), .B2(n443), .C1(n2048), .C2(n444), .A(n445), 
        .ZN(n430) );
  OAI22_X1 U488 ( .A1(n898), .A2(n102), .B1(n930), .B2(n2051), .ZN(n445) );
  OAI22_X1 U489 ( .A1(n1023), .A2(n2137), .B1(n1055), .B2(n2146), .ZN(n356) );
  OAI22_X1 U490 ( .A1(n1034), .A2(n2136), .B1(n1066), .B2(n2146), .ZN(n692) );
  OAI22_X1 U491 ( .A1(n1010), .A2(n2139), .B1(n1042), .B2(n2146), .ZN(n260) );
  OAI22_X1 U492 ( .A1(n1035), .A2(n2136), .B1(n1067), .B2(n2146), .ZN(n212) );
  OAI22_X1 U493 ( .A1(n1038), .A2(n2142), .B1(n1070), .B2(n2146), .ZN(n308) );
  OAI22_X1 U494 ( .A1(n1014), .A2(n2145), .B1(n1046), .B2(n2146), .ZN(n644) );
  OAI22_X1 U495 ( .A1(n1031), .A2(n2142), .B1(n1063), .B2(n2146), .ZN(n596) );
  OAI22_X1 U496 ( .A1(n1028), .A2(n2139), .B1(n1060), .B2(n2146), .ZN(n500) );
  OAI22_X1 U497 ( .A1(n1017), .A2(n2138), .B1(n1049), .B2(n2146), .ZN(n548) );
  OAI22_X1 U498 ( .A1(n1025), .A2(n2145), .B1(n1057), .B2(n2146), .ZN(n404) );
  OAI22_X1 U499 ( .A1(n1020), .A2(n2136), .B1(n1052), .B2(n2146), .ZN(n452) );
  OAI22_X1 U500 ( .A1(n831), .A2(n2077), .B1(n863), .B2(n2079), .ZN(n362) );
  OAI22_X1 U501 ( .A1(n842), .A2(n2077), .B1(n874), .B2(n2079), .ZN(n705) );
  OAI22_X1 U502 ( .A1(n818), .A2(n2077), .B1(n850), .B2(n2079), .ZN(n266) );
  OAI22_X1 U503 ( .A1(n843), .A2(n2077), .B1(n875), .B2(n2079), .ZN(n218) );
  OAI22_X1 U504 ( .A1(n846), .A2(n2077), .B1(n878), .B2(n2079), .ZN(n314) );
  OAI22_X1 U505 ( .A1(n822), .A2(n2077), .B1(n854), .B2(n2079), .ZN(n650) );
  OAI22_X1 U506 ( .A1(n839), .A2(n2077), .B1(n871), .B2(n2079), .ZN(n602) );
  OAI22_X1 U507 ( .A1(n836), .A2(n2077), .B1(n868), .B2(n2079), .ZN(n506) );
  OAI22_X1 U508 ( .A1(n825), .A2(n2077), .B1(n857), .B2(n2079), .ZN(n554) );
  OAI22_X1 U509 ( .A1(n828), .A2(n2077), .B1(n860), .B2(n2079), .ZN(n458) );
  OAI22_X1 U510 ( .A1(n1012), .A2(n2135), .B1(n1044), .B2(n117), .ZN(n196) );
  OAI22_X1 U511 ( .A1(n1013), .A2(n2135), .B1(n1045), .B2(n117), .ZN(n676) );
  OAI22_X1 U512 ( .A1(n1033), .A2(n2134), .B1(n1065), .B2(n2147), .ZN(n660) );
  OAI22_X1 U513 ( .A1(n1036), .A2(n2138), .B1(n1068), .B2(n117), .ZN(n244) );
  OAI22_X1 U514 ( .A1(n1011), .A2(n2137), .B1(n1043), .B2(n2147), .ZN(n228) );
  OAI22_X1 U515 ( .A1(n1008), .A2(n2140), .B1(n1040), .B2(n2147), .ZN(n324) );
  OAI22_X1 U516 ( .A1(n1009), .A2(n2141), .B1(n1041), .B2(n117), .ZN(n292) );
  OAI22_X1 U517 ( .A1(n1037), .A2(n2140), .B1(n1069), .B2(n2147), .ZN(n276) );
  OAI22_X1 U518 ( .A1(n1032), .A2(n2144), .B1(n1064), .B2(n117), .ZN(n628) );
  OAI22_X1 U519 ( .A1(n1015), .A2(n2143), .B1(n1047), .B2(n2147), .ZN(n612) );
  OAI22_X1 U520 ( .A1(n1018), .A2(n2142), .B1(n1050), .B2(n2147), .ZN(n516) );
  OAI22_X1 U521 ( .A1(n1019), .A2(n2138), .B1(n1051), .B2(n117), .ZN(n484) );
  OAI22_X1 U522 ( .A1(n1027), .A2(n2137), .B1(n1059), .B2(n2147), .ZN(n468) );
  OAI22_X1 U523 ( .A1(n1016), .A2(n2141), .B1(n1048), .B2(n117), .ZN(n580) );
  OAI22_X1 U524 ( .A1(n1030), .A2(n2140), .B1(n1062), .B2(n2147), .ZN(n564) );
  OAI22_X1 U525 ( .A1(n1029), .A2(n2143), .B1(n1061), .B2(n117), .ZN(n532) );
  OAI22_X1 U526 ( .A1(n1024), .A2(n2143), .B1(n1056), .B2(n2147), .ZN(n372) );
  OAI22_X1 U527 ( .A1(n1039), .A2(n2141), .B1(n1071), .B2(n117), .ZN(n340) );
  OAI22_X1 U528 ( .A1(n1021), .A2(n2134), .B1(n1053), .B2(n2147), .ZN(n420) );
  OAI22_X1 U529 ( .A1(n820), .A2(n95), .B1(n852), .B2(n99), .ZN(n202) );
  OAI22_X1 U530 ( .A1(n821), .A2(n95), .B1(n853), .B2(n99), .ZN(n682) );
  OAI22_X1 U531 ( .A1(n841), .A2(n2078), .B1(n873), .B2(n2080), .ZN(n666) );
  OAI22_X1 U532 ( .A1(n844), .A2(n95), .B1(n876), .B2(n99), .ZN(n250) );
  OAI22_X1 U533 ( .A1(n819), .A2(n2078), .B1(n851), .B2(n2080), .ZN(n234) );
  OAI22_X1 U534 ( .A1(n816), .A2(n2078), .B1(n848), .B2(n2080), .ZN(n330) );
  OAI22_X1 U535 ( .A1(n817), .A2(n95), .B1(n849), .B2(n99), .ZN(n298) );
  OAI22_X1 U536 ( .A1(n845), .A2(n2078), .B1(n877), .B2(n2080), .ZN(n282) );
  OAI22_X1 U537 ( .A1(n840), .A2(n95), .B1(n872), .B2(n99), .ZN(n634) );
  OAI22_X1 U538 ( .A1(n823), .A2(n2078), .B1(n855), .B2(n2080), .ZN(n618) );
  OAI22_X1 U539 ( .A1(n826), .A2(n2078), .B1(n858), .B2(n2080), .ZN(n522) );
  OAI22_X1 U540 ( .A1(n827), .A2(n95), .B1(n859), .B2(n99), .ZN(n490) );
  OAI22_X1 U541 ( .A1(n835), .A2(n2078), .B1(n867), .B2(n2080), .ZN(n474) );
  OAI22_X1 U542 ( .A1(n824), .A2(n95), .B1(n856), .B2(n99), .ZN(n586) );
  OAI22_X1 U543 ( .A1(n838), .A2(n2078), .B1(n870), .B2(n2080), .ZN(n570) );
  OAI22_X1 U544 ( .A1(n837), .A2(n95), .B1(n869), .B2(n99), .ZN(n538) );
  OAI22_X1 U545 ( .A1(n832), .A2(n2078), .B1(n864), .B2(n2080), .ZN(n378) );
  OAI22_X1 U546 ( .A1(n847), .A2(n95), .B1(n879), .B2(n99), .ZN(n346) );
  OAI22_X1 U547 ( .A1(n829), .A2(n2078), .B1(n861), .B2(n2080), .ZN(n426) );
  OAI22_X1 U548 ( .A1(n834), .A2(n95), .B1(n866), .B2(n99), .ZN(n442) );
  OAI22_X1 U549 ( .A1(n906), .A2(n2049), .B1(n938), .B2(n2051), .ZN(n710) );
  OAI22_X1 U550 ( .A1(n885), .A2(n102), .B1(n917), .B2(n2055), .ZN(n685) );
  OAI22_X1 U551 ( .A1(n905), .A2(n2050), .B1(n937), .B2(n2054), .ZN(n669) );
  OAI22_X1 U552 ( .A1(n908), .A2(n102), .B1(n940), .B2(n2052), .ZN(n253) );
  OAI22_X1 U553 ( .A1(n883), .A2(n2050), .B1(n915), .B2(n2054), .ZN(n237) );
  OAI22_X1 U554 ( .A1(n907), .A2(n2049), .B1(n939), .B2(n2053), .ZN(n221) );
  OAI22_X1 U555 ( .A1(n910), .A2(n2049), .B1(n942), .B2(n2055), .ZN(n317) );
  OAI22_X1 U556 ( .A1(n881), .A2(n102), .B1(n913), .B2(n2051), .ZN(n301) );
  OAI22_X1 U557 ( .A1(n909), .A2(n2050), .B1(n941), .B2(n2055), .ZN(n285) );
  OAI22_X1 U558 ( .A1(n886), .A2(n2049), .B1(n918), .B2(n2052), .ZN(n653) );
  OAI22_X1 U559 ( .A1(n887), .A2(n2050), .B1(n919), .B2(n2053), .ZN(n621) );
  OAI22_X1 U560 ( .A1(n903), .A2(n2049), .B1(n935), .B2(n2052), .ZN(n605) );
  OAI22_X1 U561 ( .A1(n900), .A2(n2049), .B1(n932), .B2(n2053), .ZN(n509) );
  OAI22_X1 U562 ( .A1(n891), .A2(n102), .B1(n923), .B2(n2055), .ZN(n493) );
  OAI22_X1 U563 ( .A1(n899), .A2(n2050), .B1(n931), .B2(n2052), .ZN(n477) );
  OAI22_X1 U564 ( .A1(n902), .A2(n2050), .B1(n934), .B2(n2051), .ZN(n573) );
  OAI22_X1 U565 ( .A1(n889), .A2(n2049), .B1(n921), .B2(n2053), .ZN(n557) );
  OAI22_X1 U566 ( .A1(n901), .A2(n102), .B1(n933), .B2(n2055), .ZN(n541) );
  OAI22_X1 U567 ( .A1(n896), .A2(n2050), .B1(n928), .B2(n2054), .ZN(n381) );
  OAI22_X1 U568 ( .A1(n911), .A2(n102), .B1(n943), .B2(n2052), .ZN(n349) );
  OAI22_X1 U569 ( .A1(n74), .A2(n2173), .B1(n960), .B2(n2019), .ZN(n1573) );
  OAI22_X1 U570 ( .A1(n74), .A2(n2162), .B1(n1088), .B2(n2012), .ZN(n1701) );
  OAI22_X1 U571 ( .A1(n74), .A2(n2150), .B1(n1248), .B2(n1998), .ZN(n1861) );
  OAI22_X1 U572 ( .A1(n74), .A2(n2170), .B1(n992), .B2(n110), .ZN(n1605) );
  OAI22_X1 U573 ( .A1(n74), .A2(n2160), .B1(n1120), .B2(n2009), .ZN(n1733) );
  OAI22_X1 U574 ( .A1(n74), .A2(n2153), .B1(n1216), .B2(n2001), .ZN(n1829) );
  OAI22_X1 U575 ( .A1(n74), .A2(n2189), .B1(n800), .B2(n2194), .ZN(n1413) );
  OAI22_X1 U576 ( .A1(n74), .A2(n2004), .B1(n1184), .B2(n2154), .ZN(n1797) );
  OAI22_X1 U577 ( .A1(n74), .A2(n2014), .B1(n1056), .B2(n2164), .ZN(n1669) );
  OAI22_X1 U578 ( .A1(n74), .A2(n2026), .B1(n832), .B2(n2185), .ZN(n1445) );
  OAI22_X1 U579 ( .A1(n74), .A2(n2024), .B1(n896), .B2(n2179), .ZN(n1509) );
  OAI22_X1 U580 ( .A1(n74), .A2(n2025), .B1(n864), .B2(n2182), .ZN(n1477) );
  OAI22_X1 U581 ( .A1(n74), .A2(n2022), .B1(n928), .B2(n2178), .ZN(n1541) );
  OAI22_X1 U582 ( .A1(n74), .A2(n112), .B1(n1024), .B2(n2169), .ZN(n1637) );
  OAI22_X1 U583 ( .A1(n74), .A2(n2006), .B1(n1152), .B2(n2159), .ZN(n1765) );
  OAI22_X1 U584 ( .A1(n2199), .A2(n74), .B1(n768), .B2(n2202), .ZN(n1381) );
  OAI22_X1 U585 ( .A1(n716), .A2(n8), .B1(n2327), .B2(n10), .ZN(n1265) );
  OAI22_X1 U586 ( .A1(n717), .A2(n11), .B1(n2327), .B2(n12), .ZN(n1266) );
  OAI22_X1 U587 ( .A1(n718), .A2(n13), .B1(n2327), .B2(n14), .ZN(n1267) );
  OAI22_X1 U588 ( .A1(n719), .A2(n15), .B1(n2327), .B2(n16), .ZN(n1268) );
  OAI22_X1 U589 ( .A1(n720), .A2(n17), .B1(n2327), .B2(n18), .ZN(n1269) );
  OAI22_X1 U590 ( .A1(n721), .A2(n19), .B1(n2327), .B2(n20), .ZN(n1270) );
  OAI22_X1 U591 ( .A1(n722), .A2(n21), .B1(n2327), .B2(n22), .ZN(n1271) );
  OAI22_X1 U592 ( .A1(n723), .A2(n23), .B1(n2327), .B2(n24), .ZN(n1272) );
  OAI22_X1 U593 ( .A1(n724), .A2(n25), .B1(n2327), .B2(n26), .ZN(n1273) );
  OAI22_X1 U594 ( .A1(n725), .A2(n27), .B1(n2327), .B2(n28), .ZN(n1274) );
  OAI22_X1 U595 ( .A1(n726), .A2(n29), .B1(n2327), .B2(n30), .ZN(n1275) );
  OAI22_X1 U596 ( .A1(n727), .A2(n31), .B1(n2327), .B2(n32), .ZN(n1276) );
  OAI22_X1 U597 ( .A1(n728), .A2(n33), .B1(n2327), .B2(n34), .ZN(n1277) );
  OAI22_X1 U598 ( .A1(n729), .A2(n35), .B1(n2327), .B2(n36), .ZN(n1278) );
  OAI22_X1 U599 ( .A1(n730), .A2(n37), .B1(n2327), .B2(n38), .ZN(n1279) );
  OAI22_X1 U600 ( .A1(n731), .A2(n39), .B1(n2327), .B2(n40), .ZN(n1280) );
  OAI22_X1 U601 ( .A1(n732), .A2(n11), .B1(n12), .B2(n2328), .ZN(n1281) );
  OAI22_X1 U602 ( .A1(n733), .A2(n13), .B1(n14), .B2(n2328), .ZN(n1282) );
  OAI22_X1 U603 ( .A1(n734), .A2(n15), .B1(n16), .B2(n2328), .ZN(n1283) );
  OAI22_X1 U604 ( .A1(n735), .A2(n17), .B1(n18), .B2(n2328), .ZN(n1284) );
  OAI22_X1 U605 ( .A1(n736), .A2(n19), .B1(n20), .B2(n2328), .ZN(n1285) );
  OAI22_X1 U606 ( .A1(n737), .A2(n21), .B1(n22), .B2(n2328), .ZN(n1286) );
  OAI22_X1 U607 ( .A1(n738), .A2(n23), .B1(n24), .B2(n2328), .ZN(n1287) );
  OAI22_X1 U608 ( .A1(n739), .A2(n25), .B1(n26), .B2(n2328), .ZN(n1288) );
  OAI22_X1 U609 ( .A1(n740), .A2(n27), .B1(n28), .B2(n2328), .ZN(n1289) );
  OAI22_X1 U610 ( .A1(n741), .A2(n29), .B1(n30), .B2(n2328), .ZN(n1290) );
  OAI22_X1 U611 ( .A1(n742), .A2(n31), .B1(n32), .B2(n2328), .ZN(n1291) );
  OAI22_X1 U612 ( .A1(n743), .A2(n33), .B1(n34), .B2(n2328), .ZN(n1292) );
  OAI22_X1 U613 ( .A1(n744), .A2(n35), .B1(n36), .B2(n2328), .ZN(n1293) );
  OAI22_X1 U614 ( .A1(n745), .A2(n37), .B1(n38), .B2(n2328), .ZN(n1294) );
  OAI22_X1 U615 ( .A1(n746), .A2(n39), .B1(n40), .B2(n2328), .ZN(n1295) );
  OAI22_X1 U616 ( .A1(n752), .A2(n8), .B1(n10), .B2(n2328), .ZN(n1360) );
  OAI22_X1 U617 ( .A1(n90), .A2(n2173), .B1(n959), .B2(n2019), .ZN(n1572) );
  OAI22_X1 U618 ( .A1(n90), .A2(n2163), .B1(n1087), .B2(n2012), .ZN(n1700) );
  OAI22_X1 U619 ( .A1(n68), .A2(n2172), .B1(n951), .B2(n2019), .ZN(n1564) );
  OAI22_X1 U620 ( .A1(n69), .A2(n2173), .B1(n952), .B2(n2019), .ZN(n1565) );
  OAI22_X1 U621 ( .A1(n70), .A2(n2174), .B1(n953), .B2(n2019), .ZN(n1566) );
  OAI22_X1 U622 ( .A1(n71), .A2(n2172), .B1(n954), .B2(n2019), .ZN(n1567) );
  OAI22_X1 U623 ( .A1(n72), .A2(n2173), .B1(n955), .B2(n2019), .ZN(n1568) );
  OAI22_X1 U624 ( .A1(n73), .A2(n2174), .B1(n956), .B2(n2019), .ZN(n1569) );
  OAI22_X1 U625 ( .A1(n75), .A2(n2174), .B1(n963), .B2(n2019), .ZN(n1576) );
  OAI22_X1 U626 ( .A1(n76), .A2(n2172), .B1(n964), .B2(n2019), .ZN(n1577) );
  OAI22_X1 U627 ( .A1(n79), .A2(n2172), .B1(n967), .B2(n2019), .ZN(n1580) );
  OAI22_X1 U628 ( .A1(n87), .A2(n2173), .B1(n975), .B2(n2019), .ZN(n1588) );
  OAI22_X1 U629 ( .A1(n68), .A2(n2162), .B1(n1079), .B2(n2012), .ZN(n1692) );
  OAI22_X1 U630 ( .A1(n69), .A2(n2162), .B1(n1080), .B2(n2012), .ZN(n1693) );
  OAI22_X1 U631 ( .A1(n70), .A2(n2163), .B1(n1081), .B2(n2012), .ZN(n1694) );
  OAI22_X1 U632 ( .A1(n71), .A2(n2162), .B1(n1082), .B2(n2012), .ZN(n1695) );
  OAI22_X1 U633 ( .A1(n72), .A2(n2162), .B1(n1083), .B2(n2012), .ZN(n1696) );
  OAI22_X1 U634 ( .A1(n73), .A2(n2163), .B1(n1084), .B2(n2012), .ZN(n1697) );
  OAI22_X1 U635 ( .A1(n75), .A2(n2163), .B1(n1091), .B2(n2012), .ZN(n1704) );
  OAI22_X1 U636 ( .A1(n76), .A2(n2163), .B1(n1092), .B2(n2012), .ZN(n1705) );
  OAI22_X1 U637 ( .A1(n79), .A2(n2163), .B1(n1095), .B2(n2012), .ZN(n1708) );
  OAI22_X1 U638 ( .A1(n87), .A2(n2162), .B1(n1103), .B2(n2012), .ZN(n1716) );
  OAI22_X1 U639 ( .A1(n90), .A2(n2151), .B1(n1247), .B2(n1998), .ZN(n1860) );
  OAI22_X1 U640 ( .A1(n70), .A2(n2150), .B1(n1241), .B2(n1998), .ZN(n1854) );
  OAI22_X1 U641 ( .A1(n71), .A2(n2151), .B1(n1242), .B2(n1998), .ZN(n1855) );
  OAI22_X1 U642 ( .A1(n72), .A2(n2150), .B1(n1243), .B2(n1998), .ZN(n1856) );
  OAI22_X1 U643 ( .A1(n73), .A2(n2150), .B1(n1244), .B2(n1998), .ZN(n1857) );
  OAI22_X1 U644 ( .A1(n75), .A2(n2150), .B1(n1251), .B2(n1998), .ZN(n1864) );
  OAI22_X1 U645 ( .A1(n76), .A2(n2151), .B1(n1252), .B2(n1998), .ZN(n1865) );
  OAI22_X1 U646 ( .A1(n77), .A2(n2151), .B1(n1253), .B2(n1998), .ZN(n1866) );
  OAI22_X1 U647 ( .A1(n78), .A2(n2151), .B1(n1254), .B2(n1998), .ZN(n1867) );
  OAI22_X1 U648 ( .A1(n80), .A2(n2150), .B1(n1256), .B2(n1998), .ZN(n1869) );
  OAI22_X1 U649 ( .A1(n87), .A2(n2150), .B1(n1263), .B2(n1998), .ZN(n1876) );
  OAI22_X1 U650 ( .A1(n90), .A2(n2171), .B1(n991), .B2(n110), .ZN(n1604) );
  OAI22_X1 U651 ( .A1(n90), .A2(n2161), .B1(n1119), .B2(n2009), .ZN(n1732) );
  OAI22_X1 U652 ( .A1(n90), .A2(n2153), .B1(n1215), .B2(n2001), .ZN(n1828) );
  OAI22_X1 U653 ( .A1(n69), .A2(n2170), .B1(n984), .B2(n110), .ZN(n1597) );
  OAI22_X1 U654 ( .A1(n70), .A2(n2171), .B1(n985), .B2(n110), .ZN(n1598) );
  OAI22_X1 U655 ( .A1(n71), .A2(n2170), .B1(n986), .B2(n110), .ZN(n1599) );
  OAI22_X1 U656 ( .A1(n72), .A2(n2170), .B1(n987), .B2(n110), .ZN(n1600) );
  OAI22_X1 U657 ( .A1(n73), .A2(n2170), .B1(n988), .B2(n110), .ZN(n1601) );
  OAI22_X1 U658 ( .A1(n75), .A2(n2171), .B1(n995), .B2(n2017), .ZN(n1608) );
  OAI22_X1 U659 ( .A1(n76), .A2(n2170), .B1(n996), .B2(n2016), .ZN(n1609) );
  OAI22_X1 U660 ( .A1(n78), .A2(n2171), .B1(n998), .B2(n2017), .ZN(n1611) );
  OAI22_X1 U661 ( .A1(n84), .A2(n2170), .B1(n1004), .B2(n2017), .ZN(n1617) );
  OAI22_X1 U662 ( .A1(n87), .A2(n2170), .B1(n1007), .B2(n110), .ZN(n1620) );
  OAI22_X1 U663 ( .A1(n69), .A2(n2161), .B1(n1112), .B2(n2009), .ZN(n1725) );
  OAI22_X1 U664 ( .A1(n70), .A2(n2160), .B1(n1113), .B2(n2009), .ZN(n1726) );
  OAI22_X1 U665 ( .A1(n71), .A2(n2160), .B1(n1114), .B2(n2009), .ZN(n1727) );
  OAI22_X1 U666 ( .A1(n72), .A2(n2160), .B1(n1115), .B2(n2009), .ZN(n1728) );
  OAI22_X1 U667 ( .A1(n73), .A2(n2160), .B1(n1116), .B2(n2009), .ZN(n1729) );
  OAI22_X1 U668 ( .A1(n75), .A2(n2161), .B1(n1123), .B2(n2009), .ZN(n1736) );
  OAI22_X1 U669 ( .A1(n76), .A2(n2160), .B1(n1124), .B2(n2009), .ZN(n1737) );
  OAI22_X1 U670 ( .A1(n78), .A2(n2161), .B1(n1126), .B2(n2009), .ZN(n1739) );
  OAI22_X1 U671 ( .A1(n84), .A2(n2160), .B1(n1132), .B2(n2009), .ZN(n1745) );
  OAI22_X1 U672 ( .A1(n87), .A2(n2160), .B1(n1135), .B2(n2009), .ZN(n1748) );
  OAI22_X1 U673 ( .A1(n69), .A2(n2153), .B1(n1208), .B2(n2001), .ZN(n1821) );
  OAI22_X1 U674 ( .A1(n70), .A2(n2152), .B1(n1209), .B2(n2001), .ZN(n1822) );
  OAI22_X1 U675 ( .A1(n71), .A2(n2152), .B1(n1210), .B2(n2001), .ZN(n1823) );
  OAI22_X1 U676 ( .A1(n72), .A2(n2152), .B1(n1211), .B2(n2001), .ZN(n1824) );
  OAI22_X1 U677 ( .A1(n73), .A2(n2152), .B1(n1212), .B2(n2001), .ZN(n1825) );
  OAI22_X1 U678 ( .A1(n75), .A2(n2153), .B1(n1219), .B2(n2001), .ZN(n1832) );
  OAI22_X1 U679 ( .A1(n76), .A2(n2152), .B1(n1220), .B2(n2001), .ZN(n1833) );
  OAI22_X1 U680 ( .A1(n78), .A2(n2153), .B1(n1222), .B2(n2001), .ZN(n1835) );
  OAI22_X1 U681 ( .A1(n84), .A2(n2152), .B1(n1228), .B2(n2001), .ZN(n1841) );
  OAI22_X1 U682 ( .A1(n87), .A2(n2152), .B1(n1231), .B2(n2001), .ZN(n1844) );
  OAI22_X1 U683 ( .A1(n60), .A2(n2172), .B1(n944), .B2(n2018), .ZN(n1557) );
  OAI22_X1 U684 ( .A1(n77), .A2(n2174), .B1(n965), .B2(n2018), .ZN(n1578) );
  OAI22_X1 U685 ( .A1(n78), .A2(n2172), .B1(n966), .B2(n2018), .ZN(n1579) );
  OAI22_X1 U686 ( .A1(n80), .A2(n2174), .B1(n968), .B2(n2018), .ZN(n1581) );
  OAI22_X1 U687 ( .A1(n81), .A2(n2174), .B1(n969), .B2(n2018), .ZN(n1582) );
  OAI22_X1 U688 ( .A1(n82), .A2(n2173), .B1(n970), .B2(n2018), .ZN(n1583) );
  OAI22_X1 U689 ( .A1(n83), .A2(n2172), .B1(n971), .B2(n2018), .ZN(n1584) );
  OAI22_X1 U690 ( .A1(n84), .A2(n2173), .B1(n972), .B2(n2018), .ZN(n1585) );
  OAI22_X1 U691 ( .A1(n85), .A2(n2174), .B1(n973), .B2(n2018), .ZN(n1586) );
  OAI22_X1 U692 ( .A1(n86), .A2(n2172), .B1(n974), .B2(n2018), .ZN(n1587) );
  OAI22_X1 U693 ( .A1(n60), .A2(n2163), .B1(n1072), .B2(n2011), .ZN(n1685) );
  OAI22_X1 U694 ( .A1(n77), .A2(n2163), .B1(n1093), .B2(n2011), .ZN(n1706) );
  OAI22_X1 U695 ( .A1(n78), .A2(n2162), .B1(n1094), .B2(n2011), .ZN(n1707) );
  OAI22_X1 U696 ( .A1(n80), .A2(n2163), .B1(n1096), .B2(n2011), .ZN(n1709) );
  OAI22_X1 U697 ( .A1(n81), .A2(n2163), .B1(n1097), .B2(n2011), .ZN(n1710) );
  OAI22_X1 U698 ( .A1(n82), .A2(n2162), .B1(n1098), .B2(n2011), .ZN(n1711) );
  OAI22_X1 U699 ( .A1(n83), .A2(n2163), .B1(n1099), .B2(n2011), .ZN(n1712) );
  OAI22_X1 U700 ( .A1(n84), .A2(n2162), .B1(n1100), .B2(n2011), .ZN(n1713) );
  OAI22_X1 U701 ( .A1(n85), .A2(n2163), .B1(n1101), .B2(n2011), .ZN(n1714) );
  OAI22_X1 U702 ( .A1(n86), .A2(n2163), .B1(n1102), .B2(n2011), .ZN(n1715) );
  OAI22_X1 U703 ( .A1(n60), .A2(n2170), .B1(n976), .B2(n2016), .ZN(n1589) );
  OAI22_X1 U704 ( .A1(n77), .A2(n2170), .B1(n997), .B2(n2016), .ZN(n1610) );
  OAI22_X1 U705 ( .A1(n79), .A2(n2170), .B1(n999), .B2(n2016), .ZN(n1612) );
  OAI22_X1 U706 ( .A1(n80), .A2(n2170), .B1(n1000), .B2(n2016), .ZN(n1613) );
  OAI22_X1 U707 ( .A1(n81), .A2(n2171), .B1(n1001), .B2(n2016), .ZN(n1614) );
  OAI22_X1 U708 ( .A1(n82), .A2(n2170), .B1(n1002), .B2(n2016), .ZN(n1615) );
  OAI22_X1 U709 ( .A1(n83), .A2(n2170), .B1(n1003), .B2(n2016), .ZN(n1616) );
  OAI22_X1 U710 ( .A1(n85), .A2(n2171), .B1(n1005), .B2(n2016), .ZN(n1618) );
  OAI22_X1 U711 ( .A1(n86), .A2(n2171), .B1(n1006), .B2(n2016), .ZN(n1619) );
  OAI22_X1 U712 ( .A1(n60), .A2(n2160), .B1(n1104), .B2(n2008), .ZN(n1717) );
  OAI22_X1 U713 ( .A1(n77), .A2(n2160), .B1(n1125), .B2(n2008), .ZN(n1738) );
  OAI22_X1 U714 ( .A1(n79), .A2(n2161), .B1(n1127), .B2(n2008), .ZN(n1740) );
  OAI22_X1 U715 ( .A1(n80), .A2(n2160), .B1(n1128), .B2(n2008), .ZN(n1741) );
  OAI22_X1 U716 ( .A1(n81), .A2(n2161), .B1(n1129), .B2(n2008), .ZN(n1742) );
  OAI22_X1 U717 ( .A1(n82), .A2(n2161), .B1(n1130), .B2(n2008), .ZN(n1743) );
  OAI22_X1 U718 ( .A1(n83), .A2(n2160), .B1(n1131), .B2(n2008), .ZN(n1744) );
  OAI22_X1 U719 ( .A1(n85), .A2(n2160), .B1(n1133), .B2(n2008), .ZN(n1746) );
  OAI22_X1 U720 ( .A1(n86), .A2(n2160), .B1(n1134), .B2(n2008), .ZN(n1747) );
  OAI22_X1 U721 ( .A1(n60), .A2(n2152), .B1(n1200), .B2(n2000), .ZN(n1813) );
  OAI22_X1 U722 ( .A1(n77), .A2(n2152), .B1(n1221), .B2(n2000), .ZN(n1834) );
  OAI22_X1 U723 ( .A1(n79), .A2(n2153), .B1(n1223), .B2(n2000), .ZN(n1836) );
  OAI22_X1 U724 ( .A1(n80), .A2(n2152), .B1(n1224), .B2(n2000), .ZN(n1837) );
  OAI22_X1 U725 ( .A1(n81), .A2(n2153), .B1(n1225), .B2(n2000), .ZN(n1838) );
  OAI22_X1 U726 ( .A1(n82), .A2(n2153), .B1(n1226), .B2(n2000), .ZN(n1839) );
  OAI22_X1 U727 ( .A1(n83), .A2(n2152), .B1(n1227), .B2(n2000), .ZN(n1840) );
  OAI22_X1 U728 ( .A1(n85), .A2(n2152), .B1(n1229), .B2(n2000), .ZN(n1842) );
  OAI22_X1 U729 ( .A1(n86), .A2(n2152), .B1(n1230), .B2(n2000), .ZN(n1843) );
  OAI22_X1 U730 ( .A1(n60), .A2(n2150), .B1(n1232), .B2(n1997), .ZN(n1845) );
  OAI22_X1 U731 ( .A1(n62), .A2(n2151), .B1(n1233), .B2(n1999), .ZN(n1846) );
  OAI22_X1 U732 ( .A1(n63), .A2(n2151), .B1(n1234), .B2(n1999), .ZN(n1847) );
  OAI22_X1 U733 ( .A1(n64), .A2(n2150), .B1(n1235), .B2(n1999), .ZN(n1848) );
  OAI22_X1 U734 ( .A1(n65), .A2(n2150), .B1(n1236), .B2(n1999), .ZN(n1849) );
  OAI22_X1 U735 ( .A1(n66), .A2(n2151), .B1(n1237), .B2(n1999), .ZN(n1850) );
  OAI22_X1 U736 ( .A1(n67), .A2(n2150), .B1(n1238), .B2(n1999), .ZN(n1851) );
  OAI22_X1 U737 ( .A1(n68), .A2(n2150), .B1(n1239), .B2(n1999), .ZN(n1852) );
  OAI22_X1 U738 ( .A1(n69), .A2(n2151), .B1(n1240), .B2(n1999), .ZN(n1853) );
  OAI22_X1 U739 ( .A1(n79), .A2(n2151), .B1(n1255), .B2(n1997), .ZN(n1868) );
  OAI22_X1 U740 ( .A1(n81), .A2(n2151), .B1(n1257), .B2(n1997), .ZN(n1870) );
  OAI22_X1 U741 ( .A1(n82), .A2(n2150), .B1(n1258), .B2(n1997), .ZN(n1871) );
  OAI22_X1 U742 ( .A1(n83), .A2(n2151), .B1(n1259), .B2(n1997), .ZN(n1872) );
  OAI22_X1 U743 ( .A1(n84), .A2(n2150), .B1(n1260), .B2(n1997), .ZN(n1873) );
  OAI22_X1 U744 ( .A1(n85), .A2(n2151), .B1(n1261), .B2(n1997), .ZN(n1874) );
  OAI22_X1 U745 ( .A1(n86), .A2(n2151), .B1(n1262), .B2(n1997), .ZN(n1875) );
  OAI22_X1 U746 ( .A1(n60), .A2(n115), .B1(n1040), .B2(n2166), .ZN(n1653) );
  OAI22_X1 U747 ( .A1(n69), .A2(n2014), .B1(n1048), .B2(n2166), .ZN(n1661) );
  OAI22_X1 U748 ( .A1(n71), .A2(n2014), .B1(n1050), .B2(n2166), .ZN(n1663) );
  OAI22_X1 U749 ( .A1(n72), .A2(n2014), .B1(n1051), .B2(n2166), .ZN(n1664) );
  OAI22_X1 U750 ( .A1(n76), .A2(n115), .B1(n1060), .B2(n2166), .ZN(n1673) );
  OAI22_X1 U751 ( .A1(n84), .A2(n115), .B1(n1068), .B2(n2166), .ZN(n1681) );
  OAI22_X1 U752 ( .A1(n86), .A2(n115), .B1(n1070), .B2(n2166), .ZN(n1683) );
  OAI22_X1 U753 ( .A1(n87), .A2(n2014), .B1(n1071), .B2(n2166), .ZN(n1684) );
  OAI22_X1 U754 ( .A1(n60), .A2(n93), .B1(n816), .B2(n2186), .ZN(n1429) );
  OAI22_X1 U755 ( .A1(n68), .A2(n2026), .B1(n823), .B2(n2186), .ZN(n1436) );
  OAI22_X1 U756 ( .A1(n71), .A2(n2026), .B1(n826), .B2(n2186), .ZN(n1439) );
  OAI22_X1 U757 ( .A1(n76), .A2(n93), .B1(n836), .B2(n2186), .ZN(n1449) );
  OAI22_X1 U758 ( .A1(n78), .A2(n93), .B1(n838), .B2(n2186), .ZN(n1451) );
  OAI22_X1 U759 ( .A1(n83), .A2(n93), .B1(n843), .B2(n2186), .ZN(n1456) );
  OAI22_X1 U760 ( .A1(n86), .A2(n93), .B1(n846), .B2(n2186), .ZN(n1459) );
  OAI22_X1 U761 ( .A1(n60), .A2(n100), .B1(n880), .B2(n2180), .ZN(n1493) );
  OAI22_X1 U762 ( .A1(n68), .A2(n2024), .B1(n887), .B2(n2180), .ZN(n1500) );
  OAI22_X1 U763 ( .A1(n71), .A2(n2024), .B1(n890), .B2(n2180), .ZN(n1503) );
  OAI22_X1 U764 ( .A1(n76), .A2(n100), .B1(n900), .B2(n2180), .ZN(n1513) );
  OAI22_X1 U765 ( .A1(n78), .A2(n100), .B1(n902), .B2(n2180), .ZN(n1515) );
  OAI22_X1 U766 ( .A1(n83), .A2(n100), .B1(n907), .B2(n2180), .ZN(n1520) );
  OAI22_X1 U767 ( .A1(n86), .A2(n100), .B1(n910), .B2(n2180), .ZN(n1523) );
  OAI22_X1 U768 ( .A1(n60), .A2(n97), .B1(n848), .B2(n2184), .ZN(n1461) );
  OAI22_X1 U769 ( .A1(n69), .A2(n2025), .B1(n856), .B2(n2184), .ZN(n1469) );
  OAI22_X1 U770 ( .A1(n71), .A2(n2025), .B1(n858), .B2(n2184), .ZN(n1471) );
  OAI22_X1 U771 ( .A1(n72), .A2(n2025), .B1(n859), .B2(n2184), .ZN(n1472) );
  OAI22_X1 U772 ( .A1(n76), .A2(n97), .B1(n868), .B2(n2184), .ZN(n1481) );
  OAI22_X1 U773 ( .A1(n84), .A2(n97), .B1(n876), .B2(n2184), .ZN(n1489) );
  OAI22_X1 U774 ( .A1(n86), .A2(n97), .B1(n878), .B2(n2184), .ZN(n1491) );
  OAI22_X1 U775 ( .A1(n87), .A2(n2025), .B1(n879), .B2(n2184), .ZN(n1492) );
  OAI22_X1 U776 ( .A1(n60), .A2(n2021), .B1(n912), .B2(n2177), .ZN(n1525) );
  OAI22_X1 U777 ( .A1(n69), .A2(n2022), .B1(n920), .B2(n2177), .ZN(n1533) );
  OAI22_X1 U778 ( .A1(n71), .A2(n2022), .B1(n922), .B2(n2177), .ZN(n1535) );
  OAI22_X1 U779 ( .A1(n72), .A2(n2022), .B1(n923), .B2(n2177), .ZN(n1536) );
  OAI22_X1 U780 ( .A1(n76), .A2(n2021), .B1(n932), .B2(n2177), .ZN(n1545) );
  OAI22_X1 U781 ( .A1(n84), .A2(n2021), .B1(n940), .B2(n2177), .ZN(n1553) );
  OAI22_X1 U782 ( .A1(n86), .A2(n2021), .B1(n942), .B2(n2177), .ZN(n1555) );
  OAI22_X1 U783 ( .A1(n87), .A2(n2022), .B1(n943), .B2(n2177), .ZN(n1556) );
  OAI22_X1 U784 ( .A1(n60), .A2(n2015), .B1(n1008), .B2(n2168), .ZN(n1621) );
  OAI22_X1 U785 ( .A1(n68), .A2(n112), .B1(n1015), .B2(n2168), .ZN(n1628) );
  OAI22_X1 U786 ( .A1(n71), .A2(n112), .B1(n1018), .B2(n2168), .ZN(n1631) );
  OAI22_X1 U787 ( .A1(n76), .A2(n2015), .B1(n1028), .B2(n2168), .ZN(n1641) );
  OAI22_X1 U788 ( .A1(n78), .A2(n2015), .B1(n1030), .B2(n2168), .ZN(n1643) );
  OAI22_X1 U789 ( .A1(n83), .A2(n2015), .B1(n1035), .B2(n2168), .ZN(n1648) );
  OAI22_X1 U790 ( .A1(n86), .A2(n2015), .B1(n1038), .B2(n2168), .ZN(n1651) );
  OAI22_X1 U791 ( .A1(n60), .A2(n2005), .B1(n1136), .B2(n2158), .ZN(n1749) );
  OAI22_X1 U792 ( .A1(n69), .A2(n2006), .B1(n1144), .B2(n2158), .ZN(n1757) );
  OAI22_X1 U793 ( .A1(n71), .A2(n2006), .B1(n1146), .B2(n2158), .ZN(n1759) );
  OAI22_X1 U794 ( .A1(n72), .A2(n2006), .B1(n1147), .B2(n2158), .ZN(n1760) );
  OAI22_X1 U795 ( .A1(n76), .A2(n2005), .B1(n1156), .B2(n2158), .ZN(n1769) );
  OAI22_X1 U796 ( .A1(n84), .A2(n2005), .B1(n1164), .B2(n2158), .ZN(n1777) );
  OAI22_X1 U797 ( .A1(n86), .A2(n2005), .B1(n1166), .B2(n2158), .ZN(n1779) );
  OAI22_X1 U798 ( .A1(n87), .A2(n2006), .B1(n1167), .B2(n2158), .ZN(n1780) );
  OAI22_X1 U799 ( .A1(n63), .A2(n93), .B1(n818), .B2(n2186), .ZN(n1431) );
  OAI22_X1 U800 ( .A1(n63), .A2(n100), .B1(n882), .B2(n2180), .ZN(n1495) );
  OAI22_X1 U801 ( .A1(n63), .A2(n112), .B1(n1010), .B2(n2168), .ZN(n1623) );
  OAI22_X1 U802 ( .A1(n62), .A2(n2170), .B1(n977), .B2(n2017), .ZN(n1590) );
  OAI22_X1 U803 ( .A1(n63), .A2(n2171), .B1(n978), .B2(n2017), .ZN(n1591) );
  OAI22_X1 U804 ( .A1(n64), .A2(n2170), .B1(n979), .B2(n2017), .ZN(n1592) );
  OAI22_X1 U805 ( .A1(n65), .A2(n2170), .B1(n980), .B2(n2017), .ZN(n1593) );
  OAI22_X1 U806 ( .A1(n66), .A2(n2171), .B1(n981), .B2(n2017), .ZN(n1594) );
  OAI22_X1 U807 ( .A1(n67), .A2(n2170), .B1(n982), .B2(n2017), .ZN(n1595) );
  OAI22_X1 U808 ( .A1(n68), .A2(n2171), .B1(n983), .B2(n2017), .ZN(n1596) );
  OAI22_X1 U809 ( .A1(n62), .A2(n2160), .B1(n1105), .B2(n2010), .ZN(n1718) );
  OAI22_X1 U810 ( .A1(n63), .A2(n2161), .B1(n1106), .B2(n2010), .ZN(n1719) );
  OAI22_X1 U811 ( .A1(n64), .A2(n2161), .B1(n1107), .B2(n2010), .ZN(n1720) );
  OAI22_X1 U812 ( .A1(n65), .A2(n2160), .B1(n1108), .B2(n2010), .ZN(n1721) );
  OAI22_X1 U813 ( .A1(n66), .A2(n2161), .B1(n1109), .B2(n2010), .ZN(n1722) );
  OAI22_X1 U814 ( .A1(n67), .A2(n2160), .B1(n1110), .B2(n2010), .ZN(n1723) );
  OAI22_X1 U815 ( .A1(n68), .A2(n2160), .B1(n1111), .B2(n2010), .ZN(n1724) );
  OAI22_X1 U816 ( .A1(n62), .A2(n2152), .B1(n1201), .B2(n2002), .ZN(n1814) );
  OAI22_X1 U817 ( .A1(n63), .A2(n2153), .B1(n1202), .B2(n2002), .ZN(n1815) );
  OAI22_X1 U818 ( .A1(n64), .A2(n2153), .B1(n1203), .B2(n2002), .ZN(n1816) );
  OAI22_X1 U819 ( .A1(n65), .A2(n2152), .B1(n1204), .B2(n2002), .ZN(n1817) );
  OAI22_X1 U820 ( .A1(n66), .A2(n2153), .B1(n1205), .B2(n2002), .ZN(n1818) );
  OAI22_X1 U821 ( .A1(n67), .A2(n2152), .B1(n1206), .B2(n2002), .ZN(n1819) );
  OAI22_X1 U822 ( .A1(n68), .A2(n2152), .B1(n1207), .B2(n2002), .ZN(n1820) );
  OAI22_X1 U823 ( .A1(n67), .A2(n2014), .B1(n1046), .B2(n2165), .ZN(n1659) );
  OAI22_X1 U824 ( .A1(n68), .A2(n2014), .B1(n1047), .B2(n2165), .ZN(n1660) );
  OAI22_X1 U825 ( .A1(n73), .A2(n2014), .B1(n1052), .B2(n2164), .ZN(n1665) );
  OAI22_X1 U826 ( .A1(n90), .A2(n2014), .B1(n1055), .B2(n2165), .ZN(n1668) );
  OAI22_X1 U827 ( .A1(n78), .A2(n115), .B1(n1062), .B2(n2164), .ZN(n1675) );
  OAI22_X1 U828 ( .A1(n79), .A2(n115), .B1(n1063), .B2(n2164), .ZN(n1676) );
  OAI22_X1 U829 ( .A1(n80), .A2(n115), .B1(n1064), .B2(n2164), .ZN(n1677) );
  OAI22_X1 U830 ( .A1(n81), .A2(n115), .B1(n1065), .B2(n2165), .ZN(n1678) );
  OAI22_X1 U831 ( .A1(n82), .A2(n2014), .B1(n1066), .B2(n2165), .ZN(n1679) );
  OAI22_X1 U832 ( .A1(n83), .A2(n115), .B1(n1067), .B2(n2165), .ZN(n1680) );
  OAI22_X1 U833 ( .A1(n62), .A2(n2026), .B1(n817), .B2(n2185), .ZN(n1430) );
  OAI22_X1 U834 ( .A1(n66), .A2(n2026), .B1(n821), .B2(n2187), .ZN(n1434) );
  OAI22_X1 U835 ( .A1(n70), .A2(n2026), .B1(n825), .B2(n2185), .ZN(n1438) );
  OAI22_X1 U836 ( .A1(n72), .A2(n2026), .B1(n827), .B2(n2187), .ZN(n1440) );
  OAI22_X1 U837 ( .A1(n73), .A2(n2026), .B1(n828), .B2(n2185), .ZN(n1441) );
  OAI22_X1 U838 ( .A1(n90), .A2(n2026), .B1(n831), .B2(n2187), .ZN(n1444) );
  OAI22_X1 U839 ( .A1(n77), .A2(n2026), .B1(n837), .B2(n2185), .ZN(n1450) );
  OAI22_X1 U840 ( .A1(n79), .A2(n93), .B1(n839), .B2(n2185), .ZN(n1452) );
  OAI22_X1 U841 ( .A1(n80), .A2(n2026), .B1(n840), .B2(n2187), .ZN(n1453) );
  OAI22_X1 U842 ( .A1(n81), .A2(n2026), .B1(n841), .B2(n2187), .ZN(n1454) );
  OAI22_X1 U843 ( .A1(n85), .A2(n93), .B1(n845), .B2(n2185), .ZN(n1458) );
  OAI22_X1 U844 ( .A1(n87), .A2(n2026), .B1(n847), .B2(n2187), .ZN(n1460) );
  OAI22_X1 U845 ( .A1(n62), .A2(n2024), .B1(n881), .B2(n2179), .ZN(n1494) );
  OAI22_X1 U846 ( .A1(n65), .A2(n2024), .B1(n884), .B2(n2181), .ZN(n1497) );
  OAI22_X1 U847 ( .A1(n70), .A2(n2024), .B1(n889), .B2(n2179), .ZN(n1502) );
  OAI22_X1 U848 ( .A1(n72), .A2(n2024), .B1(n891), .B2(n2181), .ZN(n1504) );
  OAI22_X1 U849 ( .A1(n73), .A2(n2024), .B1(n892), .B2(n2179), .ZN(n1505) );
  OAI22_X1 U850 ( .A1(n90), .A2(n2024), .B1(n895), .B2(n2181), .ZN(n1508) );
  OAI22_X1 U851 ( .A1(n77), .A2(n2024), .B1(n901), .B2(n2179), .ZN(n1514) );
  OAI22_X1 U852 ( .A1(n79), .A2(n100), .B1(n903), .B2(n2179), .ZN(n1516) );
  OAI22_X1 U853 ( .A1(n80), .A2(n2024), .B1(n904), .B2(n2181), .ZN(n1517) );
  OAI22_X1 U854 ( .A1(n81), .A2(n2024), .B1(n905), .B2(n2181), .ZN(n1518) );
  OAI22_X1 U855 ( .A1(n85), .A2(n100), .B1(n909), .B2(n2179), .ZN(n1522) );
  OAI22_X1 U856 ( .A1(n87), .A2(n2024), .B1(n911), .B2(n2181), .ZN(n1524) );
  OAI22_X1 U857 ( .A1(n67), .A2(n2025), .B1(n854), .B2(n2183), .ZN(n1467) );
  OAI22_X1 U858 ( .A1(n68), .A2(n2025), .B1(n855), .B2(n2183), .ZN(n1468) );
  OAI22_X1 U859 ( .A1(n73), .A2(n2025), .B1(n860), .B2(n2182), .ZN(n1473) );
  OAI22_X1 U860 ( .A1(n90), .A2(n2025), .B1(n863), .B2(n2183), .ZN(n1476) );
  OAI22_X1 U861 ( .A1(n78), .A2(n97), .B1(n870), .B2(n2182), .ZN(n1483) );
  OAI22_X1 U862 ( .A1(n79), .A2(n97), .B1(n871), .B2(n2182), .ZN(n1484) );
  OAI22_X1 U863 ( .A1(n80), .A2(n97), .B1(n872), .B2(n2182), .ZN(n1485) );
  OAI22_X1 U864 ( .A1(n81), .A2(n97), .B1(n873), .B2(n2183), .ZN(n1486) );
  OAI22_X1 U865 ( .A1(n82), .A2(n2025), .B1(n874), .B2(n2183), .ZN(n1487) );
  OAI22_X1 U866 ( .A1(n83), .A2(n97), .B1(n875), .B2(n2183), .ZN(n1488) );
  OAI22_X1 U867 ( .A1(n66), .A2(n2022), .B1(n917), .B2(n2176), .ZN(n1530) );
  OAI22_X1 U868 ( .A1(n67), .A2(n2022), .B1(n918), .B2(n2176), .ZN(n1531) );
  OAI22_X1 U869 ( .A1(n68), .A2(n2022), .B1(n919), .B2(n2176), .ZN(n1532) );
  OAI22_X1 U870 ( .A1(n73), .A2(n2022), .B1(n924), .B2(n2175), .ZN(n1537) );
  OAI22_X1 U871 ( .A1(n90), .A2(n2022), .B1(n927), .B2(n2176), .ZN(n1540) );
  OAI22_X1 U872 ( .A1(n78), .A2(n2021), .B1(n934), .B2(n2175), .ZN(n1547) );
  OAI22_X1 U873 ( .A1(n79), .A2(n2021), .B1(n935), .B2(n2175), .ZN(n1548) );
  OAI22_X1 U874 ( .A1(n80), .A2(n2021), .B1(n936), .B2(n2175), .ZN(n1549) );
  OAI22_X1 U875 ( .A1(n81), .A2(n2021), .B1(n937), .B2(n2176), .ZN(n1550) );
  OAI22_X1 U876 ( .A1(n82), .A2(n2021), .B1(n938), .B2(n2176), .ZN(n1551) );
  OAI22_X1 U877 ( .A1(n83), .A2(n2021), .B1(n939), .B2(n2176), .ZN(n1552) );
  OAI22_X1 U878 ( .A1(n62), .A2(n2015), .B1(n1009), .B2(n2167), .ZN(n1622) );
  OAI22_X1 U879 ( .A1(n66), .A2(n112), .B1(n1013), .B2(n2169), .ZN(n1626) );
  OAI22_X1 U880 ( .A1(n70), .A2(n112), .B1(n1017), .B2(n2167), .ZN(n1630) );
  OAI22_X1 U881 ( .A1(n72), .A2(n2015), .B1(n1019), .B2(n2169), .ZN(n1632) );
  OAI22_X1 U882 ( .A1(n73), .A2(n112), .B1(n1020), .B2(n2167), .ZN(n1633) );
  OAI22_X1 U883 ( .A1(n90), .A2(n2015), .B1(n1023), .B2(n2169), .ZN(n1636) );
  OAI22_X1 U884 ( .A1(n77), .A2(n2015), .B1(n1029), .B2(n2167), .ZN(n1642) );
  OAI22_X1 U885 ( .A1(n79), .A2(n2015), .B1(n1031), .B2(n2167), .ZN(n1644) );
  OAI22_X1 U886 ( .A1(n80), .A2(n2015), .B1(n1032), .B2(n2169), .ZN(n1645) );
  OAI22_X1 U887 ( .A1(n81), .A2(n2015), .B1(n1033), .B2(n2169), .ZN(n1646) );
  OAI22_X1 U888 ( .A1(n85), .A2(n2015), .B1(n1037), .B2(n2167), .ZN(n1650) );
  OAI22_X1 U889 ( .A1(n87), .A2(n112), .B1(n1039), .B2(n2169), .ZN(n1652) );
  OAI22_X1 U890 ( .A1(n67), .A2(n2006), .B1(n1142), .B2(n2157), .ZN(n1755) );
  OAI22_X1 U891 ( .A1(n68), .A2(n2006), .B1(n1143), .B2(n2157), .ZN(n1756) );
  OAI22_X1 U892 ( .A1(n73), .A2(n2006), .B1(n1148), .B2(n2156), .ZN(n1761) );
  OAI22_X1 U893 ( .A1(n90), .A2(n2006), .B1(n1151), .B2(n2157), .ZN(n1764) );
  OAI22_X1 U894 ( .A1(n78), .A2(n2005), .B1(n1158), .B2(n2156), .ZN(n1771) );
  OAI22_X1 U895 ( .A1(n79), .A2(n2005), .B1(n1159), .B2(n2156), .ZN(n1772) );
  OAI22_X1 U896 ( .A1(n80), .A2(n2005), .B1(n1160), .B2(n2156), .ZN(n1773) );
  OAI22_X1 U897 ( .A1(n81), .A2(n2005), .B1(n1161), .B2(n2157), .ZN(n1774) );
  OAI22_X1 U898 ( .A1(n82), .A2(n2005), .B1(n1162), .B2(n2157), .ZN(n1775) );
  OAI22_X1 U899 ( .A1(n83), .A2(n2005), .B1(n1163), .B2(n2157), .ZN(n1776) );
  OAI22_X1 U900 ( .A1(n64), .A2(n93), .B1(n819), .B2(n2185), .ZN(n1432) );
  OAI22_X1 U901 ( .A1(n65), .A2(n93), .B1(n820), .B2(n2187), .ZN(n1433) );
  OAI22_X1 U902 ( .A1(n64), .A2(n100), .B1(n883), .B2(n2179), .ZN(n1496) );
  OAI22_X1 U903 ( .A1(n66), .A2(n100), .B1(n885), .B2(n2181), .ZN(n1498) );
  OAI22_X1 U904 ( .A1(n64), .A2(n112), .B1(n1011), .B2(n2167), .ZN(n1624) );
  OAI22_X1 U905 ( .A1(n65), .A2(n112), .B1(n1012), .B2(n2169), .ZN(n1625) );
  OAI22_X1 U906 ( .A1(n63), .A2(n115), .B1(n1042), .B2(n2164), .ZN(n1655) );
  OAI22_X1 U907 ( .A1(n64), .A2(n115), .B1(n1043), .B2(n2164), .ZN(n1656) );
  OAI22_X1 U908 ( .A1(n65), .A2(n115), .B1(n1044), .B2(n2164), .ZN(n1657) );
  OAI22_X1 U909 ( .A1(n66), .A2(n115), .B1(n1045), .B2(n2165), .ZN(n1658) );
  OAI22_X1 U910 ( .A1(n63), .A2(n97), .B1(n850), .B2(n2182), .ZN(n1463) );
  OAI22_X1 U911 ( .A1(n64), .A2(n97), .B1(n851), .B2(n2182), .ZN(n1464) );
  OAI22_X1 U912 ( .A1(n65), .A2(n97), .B1(n852), .B2(n2182), .ZN(n1465) );
  OAI22_X1 U913 ( .A1(n66), .A2(n97), .B1(n853), .B2(n2183), .ZN(n1466) );
  OAI22_X1 U914 ( .A1(n63), .A2(n2023), .B1(n914), .B2(n2175), .ZN(n1527) );
  OAI22_X1 U915 ( .A1(n64), .A2(n2023), .B1(n915), .B2(n2175), .ZN(n1528) );
  OAI22_X1 U916 ( .A1(n65), .A2(n2023), .B1(n916), .B2(n2175), .ZN(n1529) );
  OAI22_X1 U917 ( .A1(n63), .A2(n2007), .B1(n1138), .B2(n2156), .ZN(n1751) );
  OAI22_X1 U918 ( .A1(n64), .A2(n2007), .B1(n1139), .B2(n2156), .ZN(n1752) );
  OAI22_X1 U919 ( .A1(n65), .A2(n2007), .B1(n1140), .B2(n2156), .ZN(n1753) );
  OAI22_X1 U920 ( .A1(n66), .A2(n2007), .B1(n1141), .B2(n2157), .ZN(n1754) );
  OAI22_X1 U921 ( .A1(n62), .A2(n2014), .B1(n1041), .B2(n2165), .ZN(n1654) );
  OAI22_X1 U922 ( .A1(n70), .A2(n2014), .B1(n1049), .B2(n2166), .ZN(n1662) );
  OAI22_X1 U923 ( .A1(n75), .A2(n2014), .B1(n1059), .B2(n2166), .ZN(n1672) );
  OAI22_X1 U924 ( .A1(n77), .A2(n115), .B1(n1061), .B2(n2166), .ZN(n1674) );
  OAI22_X1 U925 ( .A1(n85), .A2(n115), .B1(n1069), .B2(n2165), .ZN(n1682) );
  OAI22_X1 U926 ( .A1(n69), .A2(n2026), .B1(n824), .B2(n2187), .ZN(n1437) );
  OAI22_X1 U927 ( .A1(n75), .A2(n2026), .B1(n835), .B2(n2186), .ZN(n1448) );
  OAI22_X1 U928 ( .A1(n82), .A2(n93), .B1(n842), .B2(n2186), .ZN(n1455) );
  OAI22_X1 U929 ( .A1(n84), .A2(n93), .B1(n844), .B2(n2186), .ZN(n1457) );
  OAI22_X1 U930 ( .A1(n69), .A2(n2024), .B1(n888), .B2(n2181), .ZN(n1501) );
  OAI22_X1 U931 ( .A1(n75), .A2(n2024), .B1(n899), .B2(n2180), .ZN(n1512) );
  OAI22_X1 U932 ( .A1(n82), .A2(n100), .B1(n906), .B2(n2180), .ZN(n1519) );
  OAI22_X1 U933 ( .A1(n84), .A2(n100), .B1(n908), .B2(n2180), .ZN(n1521) );
  OAI22_X1 U934 ( .A1(n62), .A2(n2025), .B1(n849), .B2(n2183), .ZN(n1462) );
  OAI22_X1 U935 ( .A1(n70), .A2(n2025), .B1(n857), .B2(n2184), .ZN(n1470) );
  OAI22_X1 U936 ( .A1(n75), .A2(n2025), .B1(n867), .B2(n2184), .ZN(n1480) );
  OAI22_X1 U937 ( .A1(n77), .A2(n97), .B1(n869), .B2(n2184), .ZN(n1482) );
  OAI22_X1 U938 ( .A1(n85), .A2(n97), .B1(n877), .B2(n2183), .ZN(n1490) );
  OAI22_X1 U939 ( .A1(n70), .A2(n2022), .B1(n921), .B2(n2178), .ZN(n1534) );
  OAI22_X1 U940 ( .A1(n75), .A2(n2022), .B1(n931), .B2(n2178), .ZN(n1544) );
  OAI22_X1 U941 ( .A1(n77), .A2(n2021), .B1(n933), .B2(n2178), .ZN(n1546) );
  OAI22_X1 U942 ( .A1(n85), .A2(n2021), .B1(n941), .B2(n2178), .ZN(n1554) );
  OAI22_X1 U943 ( .A1(n69), .A2(n112), .B1(n1016), .B2(n2168), .ZN(n1629) );
  OAI22_X1 U944 ( .A1(n75), .A2(n112), .B1(n1027), .B2(n2168), .ZN(n1640) );
  OAI22_X1 U945 ( .A1(n82), .A2(n2015), .B1(n1034), .B2(n2168), .ZN(n1647) );
  OAI22_X1 U946 ( .A1(n84), .A2(n2015), .B1(n1036), .B2(n2169), .ZN(n1649) );
  OAI22_X1 U947 ( .A1(n62), .A2(n2006), .B1(n1137), .B2(n2159), .ZN(n1750) );
  OAI22_X1 U948 ( .A1(n70), .A2(n2006), .B1(n1145), .B2(n2159), .ZN(n1758) );
  OAI22_X1 U949 ( .A1(n75), .A2(n2006), .B1(n1155), .B2(n2159), .ZN(n1768) );
  OAI22_X1 U950 ( .A1(n77), .A2(n2005), .B1(n1157), .B2(n2159), .ZN(n1770) );
  OAI22_X1 U951 ( .A1(n85), .A2(n2005), .B1(n1165), .B2(n2159), .ZN(n1778) );
  OAI22_X1 U952 ( .A1(n67), .A2(n93), .B1(n822), .B2(n2187), .ZN(n1435) );
  OAI22_X1 U953 ( .A1(n67), .A2(n100), .B1(n886), .B2(n2181), .ZN(n1499) );
  OAI22_X1 U954 ( .A1(n67), .A2(n112), .B1(n1014), .B2(n2167), .ZN(n1627) );
  OAI22_X1 U955 ( .A1(n62), .A2(n2023), .B1(n913), .B2(n2178), .ZN(n1526) );
  OAI22_X1 U956 ( .A1(n62), .A2(n2174), .B1(n945), .B2(n2020), .ZN(n1558) );
  OAI22_X1 U957 ( .A1(n63), .A2(n2172), .B1(n946), .B2(n2020), .ZN(n1559) );
  OAI22_X1 U958 ( .A1(n64), .A2(n2172), .B1(n947), .B2(n2020), .ZN(n1560) );
  OAI22_X1 U959 ( .A1(n65), .A2(n2173), .B1(n948), .B2(n2020), .ZN(n1561) );
  OAI22_X1 U960 ( .A1(n66), .A2(n2174), .B1(n949), .B2(n2020), .ZN(n1562) );
  OAI22_X1 U961 ( .A1(n67), .A2(n2173), .B1(n950), .B2(n2020), .ZN(n1563) );
  OAI22_X1 U962 ( .A1(n62), .A2(n2163), .B1(n1073), .B2(n2013), .ZN(n1686) );
  OAI22_X1 U963 ( .A1(n63), .A2(n2162), .B1(n1074), .B2(n2013), .ZN(n1687) );
  OAI22_X1 U964 ( .A1(n64), .A2(n2163), .B1(n1075), .B2(n2013), .ZN(n1688) );
  OAI22_X1 U965 ( .A1(n65), .A2(n2163), .B1(n1076), .B2(n2013), .ZN(n1689) );
  OAI22_X1 U966 ( .A1(n66), .A2(n2163), .B1(n1077), .B2(n2013), .ZN(n1690) );
  OAI22_X1 U967 ( .A1(n67), .A2(n2162), .B1(n1078), .B2(n2013), .ZN(n1691) );
  OAI22_X1 U968 ( .A1(n60), .A2(n2188), .B1(n784), .B2(n2197), .ZN(n1397) );
  OAI22_X1 U969 ( .A1(n62), .A2(n2189), .B1(n785), .B2(n2193), .ZN(n1398) );
  OAI22_X1 U970 ( .A1(n65), .A2(n2189), .B1(n788), .B2(n2192), .ZN(n1401) );
  OAI22_X1 U971 ( .A1(n67), .A2(n2189), .B1(n790), .B2(n2196), .ZN(n1403) );
  OAI22_X1 U972 ( .A1(n68), .A2(n2189), .B1(n791), .B2(n2196), .ZN(n1404) );
  OAI22_X1 U973 ( .A1(n69), .A2(n2189), .B1(n792), .B2(n2196), .ZN(n1405) );
  OAI22_X1 U974 ( .A1(n70), .A2(n2189), .B1(n793), .B2(n2195), .ZN(n1406) );
  OAI22_X1 U975 ( .A1(n71), .A2(n2189), .B1(n794), .B2(n2195), .ZN(n1407) );
  OAI22_X1 U976 ( .A1(n72), .A2(n2189), .B1(n795), .B2(n2195), .ZN(n1408) );
  OAI22_X1 U977 ( .A1(n73), .A2(n2189), .B1(n796), .B2(n2195), .ZN(n1409) );
  OAI22_X1 U978 ( .A1(n75), .A2(n2189), .B1(n803), .B2(n2193), .ZN(n1416) );
  OAI22_X1 U979 ( .A1(n76), .A2(n2188), .B1(n804), .B2(n2193), .ZN(n1417) );
  OAI22_X1 U980 ( .A1(n77), .A2(n2188), .B1(n805), .B2(n2193), .ZN(n1418) );
  OAI22_X1 U981 ( .A1(n78), .A2(n2188), .B1(n806), .B2(n2194), .ZN(n1419) );
  OAI22_X1 U982 ( .A1(n79), .A2(n2188), .B1(n807), .B2(n2192), .ZN(n1420) );
  OAI22_X1 U983 ( .A1(n80), .A2(n2188), .B1(n808), .B2(n2192), .ZN(n1421) );
  OAI22_X1 U984 ( .A1(n81), .A2(n2188), .B1(n809), .B2(n2192), .ZN(n1422) );
  OAI22_X1 U985 ( .A1(n82), .A2(n2188), .B1(n810), .B2(n2192), .ZN(n1423) );
  OAI22_X1 U986 ( .A1(n83), .A2(n2188), .B1(n811), .B2(n2191), .ZN(n1424) );
  OAI22_X1 U987 ( .A1(n84), .A2(n2188), .B1(n812), .B2(n2193), .ZN(n1425) );
  OAI22_X1 U988 ( .A1(n85), .A2(n2188), .B1(n813), .B2(n2191), .ZN(n1426) );
  OAI22_X1 U989 ( .A1(n86), .A2(n2188), .B1(n814), .B2(n2191), .ZN(n1427) );
  OAI22_X1 U990 ( .A1(n87), .A2(n2189), .B1(n815), .B2(n2194), .ZN(n1428) );
  OAI22_X1 U991 ( .A1(n63), .A2(n2190), .B1(n786), .B2(n2194), .ZN(n1399) );
  OAI22_X1 U992 ( .A1(n64), .A2(n2190), .B1(n787), .B2(n2196), .ZN(n1400) );
  OAI22_X1 U993 ( .A1(n66), .A2(n2190), .B1(n789), .B2(n2196), .ZN(n1402) );
  OAI22_X1 U994 ( .A1(n2200), .A2(n63), .B1(n755), .B2(n2202), .ZN(n1368) );
  OAI22_X1 U995 ( .A1(n2200), .A2(n64), .B1(n756), .B2(n2202), .ZN(n1369) );
  OAI22_X1 U996 ( .A1(n2200), .A2(n66), .B1(n758), .B2(n2201), .ZN(n1371) );
  OAI22_X1 U997 ( .A1(n2200), .A2(n67), .B1(n759), .B2(n2201), .ZN(n1372) );
  OAI22_X1 U998 ( .A1(n2190), .A2(n90), .B1(n799), .B2(n2194), .ZN(n1412) );
  OAI22_X1 U999 ( .A1(n2198), .A2(n60), .B1(n753), .B2(n2202), .ZN(n1366) );
  OAI22_X1 U1000 ( .A1(n2199), .A2(n62), .B1(n754), .B2(n2202), .ZN(n1367) );
  OAI22_X1 U1001 ( .A1(n2199), .A2(n65), .B1(n757), .B2(n2201), .ZN(n1370) );
  OAI22_X1 U1002 ( .A1(n2199), .A2(n68), .B1(n760), .B2(n2201), .ZN(n1373) );
  OAI22_X1 U1003 ( .A1(n2199), .A2(n69), .B1(n761), .B2(n2201), .ZN(n1374) );
  OAI22_X1 U1004 ( .A1(n2199), .A2(n70), .B1(n762), .B2(n2201), .ZN(n1375) );
  OAI22_X1 U1005 ( .A1(n2199), .A2(n71), .B1(n763), .B2(n2201), .ZN(n1376) );
  OAI22_X1 U1006 ( .A1(n2199), .A2(n72), .B1(n764), .B2(n2203), .ZN(n1377) );
  OAI22_X1 U1007 ( .A1(n2199), .A2(n73), .B1(n765), .B2(n2202), .ZN(n1378) );
  OAI22_X1 U1008 ( .A1(n2199), .A2(n75), .B1(n771), .B2(n2202), .ZN(n1384) );
  OAI22_X1 U1009 ( .A1(n2199), .A2(n76), .B1(n772), .B2(n2202), .ZN(n1385) );
  OAI22_X1 U1010 ( .A1(n2198), .A2(n77), .B1(n773), .B2(n2201), .ZN(n1386) );
  OAI22_X1 U1011 ( .A1(n2198), .A2(n78), .B1(n774), .B2(n2201), .ZN(n1387) );
  OAI22_X1 U1012 ( .A1(n2198), .A2(n79), .B1(n775), .B2(n2201), .ZN(n1388) );
  OAI22_X1 U1013 ( .A1(n2198), .A2(n80), .B1(n776), .B2(n2201), .ZN(n1389) );
  OAI22_X1 U1014 ( .A1(n2198), .A2(n81), .B1(n777), .B2(n2201), .ZN(n1390) );
  OAI22_X1 U1015 ( .A1(n2198), .A2(n82), .B1(n778), .B2(n2201), .ZN(n1391) );
  OAI22_X1 U1016 ( .A1(n2198), .A2(n83), .B1(n779), .B2(n2201), .ZN(n1392) );
  OAI22_X1 U1017 ( .A1(n2198), .A2(n84), .B1(n780), .B2(n2201), .ZN(n1393) );
  OAI22_X1 U1018 ( .A1(n2198), .A2(n85), .B1(n781), .B2(n2201), .ZN(n1394) );
  OAI22_X1 U1019 ( .A1(n2198), .A2(n86), .B1(n782), .B2(n2201), .ZN(n1395) );
  OAI22_X1 U1020 ( .A1(n2198), .A2(n87), .B1(n783), .B2(n2201), .ZN(n1396) );
  OAI22_X1 U1021 ( .A1(n2199), .A2(n90), .B1(n1264), .B2(n2201), .ZN(n1877) );
  OAI22_X1 U1022 ( .A1(n60), .A2(n2004), .B1(n1168), .B2(n2154), .ZN(n1781) );
  OAI22_X1 U1023 ( .A1(n62), .A2(n2003), .B1(n1169), .B2(n2155), .ZN(n1782) );
  OAI22_X1 U1024 ( .A1(n63), .A2(n2003), .B1(n1170), .B2(n2155), .ZN(n1783) );
  OAI22_X1 U1025 ( .A1(n64), .A2(n2003), .B1(n1171), .B2(n2155), .ZN(n1784) );
  OAI22_X1 U1026 ( .A1(n65), .A2(n2003), .B1(n1172), .B2(n2154), .ZN(n1785) );
  OAI22_X1 U1027 ( .A1(n66), .A2(n2003), .B1(n1173), .B2(n2154), .ZN(n1786) );
  OAI22_X1 U1028 ( .A1(n67), .A2(n2003), .B1(n1174), .B2(n2154), .ZN(n1787) );
  OAI22_X1 U1029 ( .A1(n68), .A2(n2003), .B1(n1175), .B2(n2154), .ZN(n1788) );
  OAI22_X1 U1030 ( .A1(n69), .A2(n2003), .B1(n1176), .B2(n2154), .ZN(n1789) );
  OAI22_X1 U1031 ( .A1(n70), .A2(n2003), .B1(n1177), .B2(n2154), .ZN(n1790) );
  OAI22_X1 U1032 ( .A1(n71), .A2(n2003), .B1(n1178), .B2(n2155), .ZN(n1791) );
  OAI22_X1 U1033 ( .A1(n72), .A2(n2003), .B1(n1179), .B2(n2155), .ZN(n1792) );
  OAI22_X1 U1034 ( .A1(n73), .A2(n2004), .B1(n1180), .B2(n2155), .ZN(n1793) );
  OAI22_X1 U1035 ( .A1(n90), .A2(n2004), .B1(n1183), .B2(n2154), .ZN(n1796) );
  OAI22_X1 U1036 ( .A1(n75), .A2(n2004), .B1(n1187), .B2(n2154), .ZN(n1800) );
  OAI22_X1 U1037 ( .A1(n76), .A2(n2004), .B1(n1188), .B2(n2154), .ZN(n1801) );
  OAI22_X1 U1038 ( .A1(n77), .A2(n2004), .B1(n1189), .B2(n2154), .ZN(n1802) );
  OAI22_X1 U1039 ( .A1(n78), .A2(n2004), .B1(n1190), .B2(n2154), .ZN(n1803) );
  OAI22_X1 U1040 ( .A1(n79), .A2(n2004), .B1(n1191), .B2(n2155), .ZN(n1804) );
  OAI22_X1 U1041 ( .A1(n80), .A2(n2004), .B1(n1192), .B2(n2155), .ZN(n1805) );
  OAI22_X1 U1042 ( .A1(n81), .A2(n2004), .B1(n1193), .B2(n2155), .ZN(n1806) );
  OAI22_X1 U1043 ( .A1(n86), .A2(n2004), .B1(n1198), .B2(n2154), .ZN(n1811) );
  OAI22_X1 U1044 ( .A1(n87), .A2(n2003), .B1(n1199), .B2(n2154), .ZN(n1812) );
  OAI22_X1 U1045 ( .A1(n82), .A2(n2004), .B1(n1194), .B2(n2154), .ZN(n1807) );
  OAI22_X1 U1046 ( .A1(n83), .A2(n127), .B1(n1195), .B2(n2154), .ZN(n1808) );
  OAI22_X1 U1047 ( .A1(n84), .A2(n2003), .B1(n1196), .B2(n2154), .ZN(n1809) );
  OAI22_X1 U1048 ( .A1(n85), .A2(n127), .B1(n1197), .B2(n2154), .ZN(n1810) );
  NAND4_X1 U1049 ( .A1(n622), .A2(n623), .A3(n624), .A4(n625), .ZN(N104) );
  AOI221_X1 U1050 ( .B1(n2060), .B2(n632), .C1(n2075), .C2(n633), .A(n634), 
        .ZN(n623) );
  AOI221_X1 U1051 ( .B1(n2115), .B2(n626), .C1(n2130), .C2(n627), .A(n628), 
        .ZN(n625) );
  NAND4_X1 U1052 ( .A1(n190), .A2(n191), .A3(n192), .A4(n193), .ZN(N99) );
  AOI221_X1 U1053 ( .B1(n2058), .B2(n200), .C1(n2066), .C2(n201), .A(n202), 
        .ZN(n191) );
  AOI221_X1 U1054 ( .B1(n2113), .B2(n194), .C1(n2121), .C2(n195), .A(n196), 
        .ZN(n193) );
  NAND4_X1 U1055 ( .A1(n254), .A2(n255), .A3(n256), .A4(n257), .ZN(N95) );
  AOI221_X1 U1056 ( .B1(n2112), .B2(n258), .C1(n2125), .C2(n259), .A(n260), 
        .ZN(n257) );
  AOI221_X1 U1057 ( .B1(n2057), .B2(n264), .C1(n2070), .C2(n265), .A(n266), 
        .ZN(n255) );
  NAND4_X1 U1058 ( .A1(n318), .A2(n319), .A3(n320), .A4(n321), .ZN(N91) );
  AOI221_X1 U1059 ( .B1(n2059), .B2(n328), .C1(n2071), .C2(n329), .A(n330), 
        .ZN(n319) );
  AOI221_X1 U1060 ( .B1(n2114), .B2(n322), .C1(n2126), .C2(n323), .A(n324), 
        .ZN(n321) );
  NAND4_X1 U1061 ( .A1(n510), .A2(n511), .A3(n512), .A4(n513), .ZN(N111) );
  AOI221_X1 U1062 ( .B1(n2057), .B2(n520), .C1(n2073), .C2(n521), .A(n522), 
        .ZN(n511) );
  AOI221_X1 U1063 ( .B1(n2112), .B2(n514), .C1(n2128), .C2(n515), .A(n516), 
        .ZN(n513) );
  NAND4_X1 U1064 ( .A1(n574), .A2(n575), .A3(n576), .A4(n577), .ZN(N107) );
  AOI221_X1 U1065 ( .B1(n2058), .B2(n584), .C1(n2072), .C2(n585), .A(n586), 
        .ZN(n575) );
  AOI221_X1 U1066 ( .B1(n2113), .B2(n578), .C1(n2127), .C2(n579), .A(n580), 
        .ZN(n577) );
  AOI221_X1 U1067 ( .B1(n2061), .B2(n424), .C1(n2065), .C2(n425), .A(n426), 
        .ZN(n415) );
  AOI221_X1 U1068 ( .B1(n2116), .B2(n418), .C1(n2120), .C2(n419), .A(n420), 
        .ZN(n417) );
  AOI221_X1 U1069 ( .B1(n2062), .B2(n440), .C1(n2066), .C2(n441), .A(n442), 
        .ZN(n431) );
  NAND4_X1 U1070 ( .A1(n382), .A2(n383), .A3(n384), .A4(n385), .ZN(N119) );
  NAND4_X1 U1071 ( .A1(n398), .A2(n399), .A3(n400), .A4(n401), .ZN(N118) );
  NAND4_X1 U1072 ( .A1(n446), .A2(n447), .A3(n448), .A4(n449), .ZN(N115) );
  AOI221_X1 U1073 ( .B1(n2114), .B2(n450), .C1(n2122), .C2(n451), .A(n452), 
        .ZN(n449) );
  AOI221_X1 U1074 ( .B1(n2059), .B2(n456), .C1(n2067), .C2(n457), .A(n458), 
        .ZN(n447) );
  OAI21_X1 U1075 ( .B1(n2235), .B2(n2228), .A(n2227), .ZN(PRED[0]) );
  NAND2_X1 U1076 ( .A1(n2200), .A2(n766), .ZN(n1379) );
  NAND2_X1 U1077 ( .A1(n2200), .A2(n767), .ZN(n1380) );
  NAND2_X1 U1078 ( .A1(n2200), .A2(n769), .ZN(n1382) );
  NAND2_X1 U1079 ( .A1(n2200), .A2(n770), .ZN(n1383) );
  INV_X1 U1080 ( .A(CURR_PC[2]), .ZN(n713) );
  NAND2_X1 U1081 ( .A1(n2190), .A2(n797), .ZN(n1410) );
  NAND2_X1 U1082 ( .A1(n2190), .A2(n801), .ZN(n1414) );
  NAND2_X1 U1083 ( .A1(n2190), .A2(n802), .ZN(n1415) );
  INV_X1 U1084 ( .A(CURR_PC[4]), .ZN(n698) );
  INV_X1 U1085 ( .A(CURR_PC[5]), .ZN(n707) );
  INV_X1 U1086 ( .A(CURR_PC[3]), .ZN(n712) );
  NAND2_X1 U1089 ( .A1(n2026), .A2(n829), .ZN(n1442) );
  NAND2_X1 U1090 ( .A1(n93), .A2(n830), .ZN(n1443) );
  NAND2_X1 U1091 ( .A1(n93), .A2(n834), .ZN(n1447) );
  NAND2_X1 U1092 ( .A1(n2024), .A2(n894), .ZN(n1507) );
  NAND2_X1 U1093 ( .A1(n100), .A2(n897), .ZN(n1510) );
  NAND2_X1 U1094 ( .A1(n100), .A2(n898), .ZN(n1511) );
  NAND2_X1 U1095 ( .A1(n2015), .A2(n1021), .ZN(n1634) );
  NAND2_X1 U1096 ( .A1(n112), .A2(n1022), .ZN(n1635) );
  NAND2_X1 U1097 ( .A1(n112), .A2(n1025), .ZN(n1638) );
  NAND2_X1 U1098 ( .A1(n2173), .A2(n958), .ZN(n1571) );
  NAND2_X1 U1099 ( .A1(n2162), .A2(n1085), .ZN(n1698) );
  NAND2_X1 U1100 ( .A1(n2174), .A2(n962), .ZN(n1575) );
  NAND2_X1 U1101 ( .A1(n2171), .A2(n994), .ZN(n1607) );
  NAND2_X1 U1102 ( .A1(n2163), .A2(n1086), .ZN(n1699) );
  NAND2_X1 U1103 ( .A1(n2161), .A2(n1117), .ZN(n1730) );
  NAND2_X1 U1104 ( .A1(n2153), .A2(n1214), .ZN(n1827) );
  NAND2_X1 U1105 ( .A1(n127), .A2(n1185), .ZN(n1798) );
  NAND2_X1 U1106 ( .A1(n2014), .A2(n1053), .ZN(n1666) );
  NAND2_X1 U1107 ( .A1(n115), .A2(n1057), .ZN(n1670) );
  NAND2_X1 U1108 ( .A1(n2025), .A2(n861), .ZN(n1474) );
  NAND2_X1 U1109 ( .A1(n97), .A2(n866), .ZN(n1479) );
  NAND2_X1 U1110 ( .A1(n2023), .A2(n929), .ZN(n1542) );
  NAND2_X1 U1111 ( .A1(n2023), .A2(n930), .ZN(n1543) );
  NAND2_X1 U1112 ( .A1(n2007), .A2(n1150), .ZN(n1763) );
  NAND2_X1 U1113 ( .A1(n2007), .A2(n1153), .ZN(n1766) );
  INV_X1 U1114 ( .A(CURR_PC[0]), .ZN(n90) );
  INV_X1 U1115 ( .A(CURR_PC[30]), .ZN(n60) );
  INV_X1 U1116 ( .A(CURR_PC[28]), .ZN(n62) );
  INV_X1 U1117 ( .A(CURR_PC[26]), .ZN(n63) );
  INV_X1 U1118 ( .A(CURR_PC[24]), .ZN(n64) );
  INV_X1 U1119 ( .A(CURR_PC[22]), .ZN(n65) );
  INV_X1 U1120 ( .A(CURR_PC[20]), .ZN(n66) );
  INV_X1 U1121 ( .A(CURR_PC[18]), .ZN(n67) );
  INV_X1 U1122 ( .A(CURR_PC[16]), .ZN(n68) );
  INV_X1 U1123 ( .A(CURR_PC[14]), .ZN(n69) );
  INV_X1 U1124 ( .A(CURR_PC[12]), .ZN(n70) );
  INV_X1 U1125 ( .A(CURR_PC[10]), .ZN(n71) );
  INV_X1 U1126 ( .A(CURR_PC[8]), .ZN(n72) );
  INV_X1 U1127 ( .A(CURR_PC[6]), .ZN(n73) );
  INV_X1 U1128 ( .A(CURR_PC[7]), .ZN(n75) );
  INV_X1 U1129 ( .A(CURR_PC[9]), .ZN(n76) );
  INV_X1 U1130 ( .A(CURR_PC[11]), .ZN(n77) );
  INV_X1 U1131 ( .A(CURR_PC[13]), .ZN(n78) );
  INV_X1 U1132 ( .A(CURR_PC[15]), .ZN(n79) );
  INV_X1 U1133 ( .A(CURR_PC[17]), .ZN(n80) );
  INV_X1 U1134 ( .A(CURR_PC[19]), .ZN(n81) );
  INV_X1 U1135 ( .A(CURR_PC[21]), .ZN(n82) );
  INV_X1 U1136 ( .A(CURR_PC[23]), .ZN(n83) );
  INV_X1 U1137 ( .A(CURR_PC[25]), .ZN(n84) );
  INV_X1 U1138 ( .A(CURR_PC[27]), .ZN(n85) );
  INV_X1 U1139 ( .A(CURR_PC[29]), .ZN(n86) );
  INV_X1 U1140 ( .A(CURR_PC[31]), .ZN(n87) );
  NOR2_X1 U1141 ( .A1(n748), .A2(n750), .ZN(n50) );
  NOR2_X1 U1142 ( .A1(\PC_HISTORY[1][2] ), .A2(n750), .ZN(n49) );
  NOR2_X1 U1143 ( .A1(\PC_HISTORY[1][3] ), .A2(n748), .ZN(n48) );
  AOI221_X1 U1144 ( .B1(n2030), .B2(\PRED_TABLE[8][1] ), .C1(n2043), .C2(
        \PRED_TABLE[9][1] ), .A(n189), .ZN(n174) );
  OAI22_X1 U1145 ( .A1(n737), .A2(n2050), .B1(n741), .B2(n2051), .ZN(n189) );
  OAI22_X1 U1146 ( .A1(n735), .A2(n2134), .B1(n743), .B2(n2147), .ZN(n180) );
  OAI22_X1 U1147 ( .A1(n738), .A2(n2078), .B1(n740), .B2(n2080), .ZN(n186) );
  OAI22_X1 U1148 ( .A1(n733), .A2(n2098), .B1(n745), .B2(n2105), .ZN(n183) );
  AND2_X1 U1149 ( .A1(n751), .A2(n57), .ZN(n53) );
  AND2_X1 U1150 ( .A1(n751), .A2(n51), .ZN(n54) );
  AND2_X1 U1152 ( .A1(n747), .A2(MISS_HIT[1]), .ZN(n51) );
  MUX2_X1 U1153 ( .A(\PRED_TABLE[7][0] ), .B(\PRED_TABLE[15][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1966) );
  MUX2_X1 U1154 ( .A(\PRED_TABLE[3][0] ), .B(\PRED_TABLE[11][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1967) );
  MUX2_X1 U1155 ( .A(n1967), .B(n1966), .S(\PC_HISTORY[1][2] ), .Z(n1968) );
  MUX2_X1 U1156 ( .A(\PRED_TABLE[6][0] ), .B(\PRED_TABLE[14][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1969) );
  MUX2_X1 U1157 ( .A(\PRED_TABLE[2][0] ), .B(\PRED_TABLE[10][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1970) );
  MUX2_X1 U1158 ( .A(n1970), .B(n1969), .S(\PC_HISTORY[1][2] ), .Z(n1971) );
  MUX2_X1 U1159 ( .A(n1971), .B(n1968), .S(\PC_HISTORY[1][0] ), .Z(n1972) );
  MUX2_X1 U1160 ( .A(\PRED_TABLE[5][0] ), .B(\PRED_TABLE[13][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1973) );
  MUX2_X1 U1161 ( .A(\PRED_TABLE[1][0] ), .B(\PRED_TABLE[9][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1974) );
  MUX2_X1 U1162 ( .A(n1974), .B(n1973), .S(\PC_HISTORY[1][2] ), .Z(n1975) );
  MUX2_X1 U1163 ( .A(\PRED_TABLE[4][0] ), .B(\PRED_TABLE[12][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1976) );
  MUX2_X1 U1164 ( .A(\PRED_TABLE[0][0] ), .B(\PRED_TABLE[8][0] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1977) );
  MUX2_X1 U1165 ( .A(n1977), .B(n1976), .S(\PC_HISTORY[1][2] ), .Z(n1978) );
  MUX2_X1 U1166 ( .A(n1978), .B(n1975), .S(\PC_HISTORY[1][0] ), .Z(n1979) );
  MUX2_X1 U1167 ( .A(n1979), .B(n1972), .S(\PC_HISTORY[1][1] ), .Z(N850) );
  MUX2_X1 U1168 ( .A(\PRED_TABLE[7][1] ), .B(\PRED_TABLE[15][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1980) );
  MUX2_X1 U1169 ( .A(\PRED_TABLE[3][1] ), .B(\PRED_TABLE[11][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1981) );
  MUX2_X1 U1170 ( .A(n1981), .B(n1980), .S(\PC_HISTORY[1][2] ), .Z(n1982) );
  MUX2_X1 U1171 ( .A(\PRED_TABLE[6][1] ), .B(\PRED_TABLE[14][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1983) );
  MUX2_X1 U1172 ( .A(\PRED_TABLE[2][1] ), .B(\PRED_TABLE[10][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1984) );
  MUX2_X1 U1173 ( .A(n1984), .B(n1983), .S(\PC_HISTORY[1][2] ), .Z(n1985) );
  MUX2_X1 U1174 ( .A(n1985), .B(n1982), .S(\PC_HISTORY[1][0] ), .Z(n1986) );
  MUX2_X1 U1175 ( .A(\PRED_TABLE[5][1] ), .B(\PRED_TABLE[13][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1987) );
  MUX2_X1 U1176 ( .A(\PRED_TABLE[1][1] ), .B(\PRED_TABLE[9][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1988) );
  MUX2_X1 U1177 ( .A(n1988), .B(n1987), .S(\PC_HISTORY[1][2] ), .Z(n1989) );
  MUX2_X1 U1178 ( .A(\PRED_TABLE[4][1] ), .B(\PRED_TABLE[12][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1990) );
  MUX2_X1 U1179 ( .A(\PRED_TABLE[0][1] ), .B(\PRED_TABLE[8][1] ), .S(
        \PC_HISTORY[1][3] ), .Z(n1991) );
  MUX2_X1 U1180 ( .A(n1991), .B(n1990), .S(\PC_HISTORY[1][2] ), .Z(n1992) );
  MUX2_X1 U1181 ( .A(n1992), .B(n1989), .S(\PC_HISTORY[1][0] ), .Z(n1993) );
  MUX2_X1 U1182 ( .A(n1993), .B(n1986), .S(\PC_HISTORY[1][1] ), .Z(N849) );
  OAI21_X1 U1183 ( .B1(n2235), .B2(n2232), .A(n2231), .ZN(PRED[1]) );
  NAND2_X1 U1184 ( .A1(n2326), .A2(n1964), .ZN(PRED[31]) );
  INV_X1 U1185 ( .A(CURR_PC[1]), .ZN(n74) );
  NAND2_X1 U1186 ( .A1(n1963), .A2(MISS_HIT[1]), .ZN(n2223) );
  INV_X1 U1187 ( .A(n2197), .ZN(n2190) );
  INV_X1 U1188 ( .A(n2203), .ZN(n2200) );
  CLKBUF_X1 U1189 ( .A(n2215), .Z(n2205) );
  CLKBUF_X1 U1190 ( .A(n2215), .Z(n2206) );
  CLKBUF_X1 U1191 ( .A(n2215), .Z(n2207) );
  CLKBUF_X1 U1192 ( .A(n2215), .Z(n2208) );
  CLKBUF_X1 U1193 ( .A(n2214), .Z(n2209) );
  CLKBUF_X1 U1194 ( .A(n2214), .Z(n2210) );
  CLKBUF_X1 U1195 ( .A(n2214), .Z(n2211) );
  CLKBUF_X1 U1196 ( .A(n2214), .Z(n2212) );
  CLKBUF_X1 U1197 ( .A(n2214), .Z(n2213) );
  INV_X1 U1199 ( .A(INST_27), .ZN(n2216) );
  NAND3_X1 U1200 ( .A1(INST_28), .A2(n715), .A3(n2216), .ZN(n2224) );
  INV_X1 U1203 ( .A(n2366), .ZN(n2329) );
  INV_X1 U1204 ( .A(N850), .ZN(n2218) );
  INV_X1 U1205 ( .A(N849), .ZN(n2220) );
  NAND4_X1 U1207 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(n2222) );
  INV_X1 U1209 ( .A(n2323), .ZN(n2235) );
  INV_X1 U1210 ( .A(NEXT_PC[0]), .ZN(n2228) );
  INV_X1 U1211 ( .A(NEW_PC[0]), .ZN(n2225) );
  AOI21_X1 U1212 ( .B1(PRED_TK[0]), .B2(n1994), .A(n2226), .ZN(n2227) );
  INV_X1 U1213 ( .A(NEXT_PC[1]), .ZN(n2232) );
  INV_X1 U1214 ( .A(NEW_PC[1]), .ZN(n2229) );
  AOI21_X1 U1215 ( .B1(PRED_TK[1]), .B2(n1994), .A(n2230), .ZN(n2231) );
  INV_X1 U1216 ( .A(NEW_PC[2]), .ZN(n2236) );
  INV_X1 U1217 ( .A(NEXT_PC[2]), .ZN(n2234) );
  NAND2_X1 U1218 ( .A1(PRED_TK[2]), .A2(n1994), .ZN(n2233) );
  NAND2_X1 U1220 ( .A1(PRED_TK[3]), .A2(n1994), .ZN(n2240) );
  NAND2_X1 U1221 ( .A1(NEW_PC[3]), .A2(n2322), .ZN(n2239) );
  NAND2_X1 U1222 ( .A1(NEXT_PC[3]), .A2(n2027), .ZN(n2238) );
  NAND3_X1 U1223 ( .A1(n2240), .A2(n2239), .A3(n2238), .ZN(PRED[3]) );
  NAND2_X1 U1224 ( .A1(PRED_TK[4]), .A2(n1994), .ZN(n2243) );
  NAND2_X1 U1225 ( .A1(NEW_PC[4]), .A2(n2322), .ZN(n2242) );
  NAND2_X1 U1226 ( .A1(NEXT_PC[4]), .A2(n2323), .ZN(n2241) );
  NAND3_X1 U1227 ( .A1(n2243), .A2(n2242), .A3(n2241), .ZN(PRED[4]) );
  NAND2_X1 U1228 ( .A1(PRED_TK[5]), .A2(n1994), .ZN(n2246) );
  NAND2_X1 U1229 ( .A1(NEW_PC[5]), .A2(n2322), .ZN(n2245) );
  NAND2_X1 U1230 ( .A1(NEXT_PC[5]), .A2(n2027), .ZN(n2244) );
  NAND3_X1 U1231 ( .A1(n2246), .A2(n2245), .A3(n2244), .ZN(PRED[5]) );
  NAND2_X1 U1232 ( .A1(PRED_TK[6]), .A2(n1994), .ZN(n2249) );
  NAND2_X1 U1233 ( .A1(NEW_PC[6]), .A2(n2322), .ZN(n2248) );
  NAND2_X1 U1234 ( .A1(NEXT_PC[6]), .A2(n2323), .ZN(n2247) );
  NAND3_X1 U1235 ( .A1(n2249), .A2(n2248), .A3(n2247), .ZN(PRED[6]) );
  NAND2_X1 U1236 ( .A1(PRED_TK[7]), .A2(n1994), .ZN(n2252) );
  NAND2_X1 U1237 ( .A1(NEW_PC[7]), .A2(n2322), .ZN(n2251) );
  NAND2_X1 U1238 ( .A1(NEXT_PC[7]), .A2(n2027), .ZN(n2250) );
  NAND3_X1 U1239 ( .A1(n2252), .A2(n2251), .A3(n2250), .ZN(PRED[7]) );
  NAND2_X1 U1240 ( .A1(PRED_TK[8]), .A2(n1994), .ZN(n2255) );
  NAND2_X1 U1241 ( .A1(NEW_PC[8]), .A2(n2322), .ZN(n2254) );
  NAND2_X1 U1242 ( .A1(NEXT_PC[8]), .A2(n2323), .ZN(n2253) );
  NAND3_X1 U1243 ( .A1(n2255), .A2(n2254), .A3(n2253), .ZN(PRED[8]) );
  NAND2_X1 U1244 ( .A1(PRED_TK[9]), .A2(n1994), .ZN(n2258) );
  NAND2_X1 U1245 ( .A1(NEW_PC[9]), .A2(n2322), .ZN(n2257) );
  NAND2_X1 U1246 ( .A1(NEXT_PC[9]), .A2(n2027), .ZN(n2256) );
  NAND3_X1 U1247 ( .A1(n2258), .A2(n2257), .A3(n2256), .ZN(PRED[9]) );
  NAND2_X1 U1248 ( .A1(PRED_TK[10]), .A2(n1994), .ZN(n2261) );
  NAND2_X1 U1249 ( .A1(NEW_PC[10]), .A2(n2322), .ZN(n2260) );
  NAND2_X1 U1250 ( .A1(NEXT_PC[10]), .A2(n2323), .ZN(n2259) );
  NAND3_X1 U1251 ( .A1(n2261), .A2(n2260), .A3(n2259), .ZN(PRED[10]) );
  NAND2_X1 U1252 ( .A1(PRED_TK[11]), .A2(n1994), .ZN(n2264) );
  NAND2_X1 U1253 ( .A1(NEW_PC[11]), .A2(n2322), .ZN(n2263) );
  NAND2_X1 U1254 ( .A1(NEXT_PC[11]), .A2(n2027), .ZN(n2262) );
  NAND3_X1 U1255 ( .A1(n2264), .A2(n2263), .A3(n2262), .ZN(PRED[11]) );
  NAND2_X1 U1256 ( .A1(PRED_TK[12]), .A2(n1995), .ZN(n2267) );
  NAND2_X1 U1257 ( .A1(NEW_PC[12]), .A2(n2322), .ZN(n2266) );
  NAND2_X1 U1258 ( .A1(NEXT_PC[12]), .A2(n2323), .ZN(n2265) );
  NAND3_X1 U1259 ( .A1(n2267), .A2(n2266), .A3(n2265), .ZN(PRED[12]) );
  NAND2_X1 U1260 ( .A1(PRED_TK[13]), .A2(n1995), .ZN(n2270) );
  NAND2_X1 U1261 ( .A1(NEW_PC[13]), .A2(n2322), .ZN(n2269) );
  NAND2_X1 U1262 ( .A1(NEXT_PC[13]), .A2(n2027), .ZN(n2268) );
  NAND3_X1 U1263 ( .A1(n2270), .A2(n2269), .A3(n2268), .ZN(PRED[13]) );
  NAND2_X1 U1264 ( .A1(PRED_TK[14]), .A2(n1995), .ZN(n2273) );
  NAND2_X1 U1265 ( .A1(NEW_PC[14]), .A2(n2322), .ZN(n2272) );
  NAND2_X1 U1266 ( .A1(NEXT_PC[14]), .A2(n2323), .ZN(n2271) );
  NAND3_X1 U1267 ( .A1(n2273), .A2(n2272), .A3(n2271), .ZN(PRED[14]) );
  NAND2_X1 U1268 ( .A1(PRED_TK[15]), .A2(n1995), .ZN(n2276) );
  NAND2_X1 U1269 ( .A1(NEW_PC[15]), .A2(n2322), .ZN(n2275) );
  NAND2_X1 U1270 ( .A1(NEXT_PC[15]), .A2(n2027), .ZN(n2274) );
  NAND3_X1 U1271 ( .A1(n2276), .A2(n2275), .A3(n2274), .ZN(PRED[15]) );
  NAND2_X1 U1272 ( .A1(PRED_TK[16]), .A2(n1995), .ZN(n2279) );
  NAND2_X1 U1273 ( .A1(NEW_PC[16]), .A2(n2322), .ZN(n2278) );
  NAND2_X1 U1274 ( .A1(NEXT_PC[16]), .A2(n2323), .ZN(n2277) );
  NAND3_X1 U1275 ( .A1(n2279), .A2(n2278), .A3(n2277), .ZN(PRED[16]) );
  NAND2_X1 U1276 ( .A1(PRED_TK[17]), .A2(n1995), .ZN(n2282) );
  NAND2_X1 U1277 ( .A1(NEW_PC[17]), .A2(n2322), .ZN(n2281) );
  NAND2_X1 U1278 ( .A1(NEXT_PC[17]), .A2(n2027), .ZN(n2280) );
  NAND3_X1 U1279 ( .A1(n2282), .A2(n2281), .A3(n2280), .ZN(PRED[17]) );
  NAND2_X1 U1280 ( .A1(PRED_TK[18]), .A2(n1995), .ZN(n2285) );
  NAND2_X1 U1281 ( .A1(NEW_PC[18]), .A2(n2322), .ZN(n2284) );
  NAND2_X1 U1282 ( .A1(NEXT_PC[18]), .A2(n2323), .ZN(n2283) );
  NAND3_X1 U1283 ( .A1(n2285), .A2(n2284), .A3(n2283), .ZN(PRED[18]) );
  NAND2_X1 U1284 ( .A1(PRED_TK[19]), .A2(n1995), .ZN(n2288) );
  NAND2_X1 U1285 ( .A1(NEW_PC[19]), .A2(n2322), .ZN(n2287) );
  NAND2_X1 U1286 ( .A1(NEXT_PC[19]), .A2(n2027), .ZN(n2286) );
  NAND3_X1 U1287 ( .A1(n2288), .A2(n2287), .A3(n2286), .ZN(PRED[19]) );
  NAND2_X1 U1288 ( .A1(PRED_TK[20]), .A2(n1995), .ZN(n2291) );
  NAND2_X1 U1289 ( .A1(NEW_PC[20]), .A2(n2322), .ZN(n2290) );
  NAND2_X1 U1290 ( .A1(NEXT_PC[20]), .A2(n2323), .ZN(n2289) );
  NAND3_X1 U1291 ( .A1(n2291), .A2(n2290), .A3(n2289), .ZN(PRED[20]) );
  NAND2_X1 U1292 ( .A1(PRED_TK[21]), .A2(n1995), .ZN(n2294) );
  NAND2_X1 U1293 ( .A1(NEW_PC[21]), .A2(n2322), .ZN(n2293) );
  NAND2_X1 U1294 ( .A1(NEXT_PC[21]), .A2(n2027), .ZN(n2292) );
  NAND3_X1 U1295 ( .A1(n2294), .A2(n2293), .A3(n2292), .ZN(PRED[21]) );
  NAND2_X1 U1296 ( .A1(PRED_TK[22]), .A2(n1995), .ZN(n2297) );
  NAND2_X1 U1297 ( .A1(NEW_PC[22]), .A2(n2322), .ZN(n2296) );
  NAND2_X1 U1298 ( .A1(NEXT_PC[22]), .A2(n2323), .ZN(n2295) );
  NAND3_X1 U1299 ( .A1(n2297), .A2(n2296), .A3(n2295), .ZN(PRED[22]) );
  NAND2_X1 U1300 ( .A1(PRED_TK[23]), .A2(n1995), .ZN(n2300) );
  NAND2_X1 U1301 ( .A1(NEW_PC[23]), .A2(n2322), .ZN(n2299) );
  NAND2_X1 U1302 ( .A1(NEXT_PC[23]), .A2(n2027), .ZN(n2298) );
  NAND3_X1 U1303 ( .A1(n2300), .A2(n2299), .A3(n2298), .ZN(PRED[23]) );
  NAND2_X1 U1304 ( .A1(PRED_TK[24]), .A2(n1996), .ZN(n2303) );
  NAND2_X1 U1305 ( .A1(NEW_PC[24]), .A2(n2322), .ZN(n2302) );
  NAND2_X1 U1306 ( .A1(NEXT_PC[24]), .A2(n2323), .ZN(n2301) );
  NAND3_X1 U1307 ( .A1(n2303), .A2(n2302), .A3(n2301), .ZN(PRED[24]) );
  NAND2_X1 U1308 ( .A1(PRED_TK[25]), .A2(n1996), .ZN(n2306) );
  NAND2_X1 U1309 ( .A1(NEW_PC[25]), .A2(n2322), .ZN(n2305) );
  NAND2_X1 U1310 ( .A1(NEXT_PC[25]), .A2(n2027), .ZN(n2304) );
  NAND3_X1 U1311 ( .A1(n2306), .A2(n2305), .A3(n2304), .ZN(PRED[25]) );
  NAND2_X1 U1312 ( .A1(PRED_TK[26]), .A2(n1996), .ZN(n2309) );
  NAND2_X1 U1313 ( .A1(NEW_PC[26]), .A2(n2322), .ZN(n2308) );
  NAND2_X1 U1314 ( .A1(NEXT_PC[26]), .A2(n2323), .ZN(n2307) );
  NAND3_X1 U1315 ( .A1(n2309), .A2(n2308), .A3(n2307), .ZN(PRED[26]) );
  NAND2_X1 U1316 ( .A1(PRED_TK[27]), .A2(n1996), .ZN(n2312) );
  NAND2_X1 U1317 ( .A1(NEW_PC[27]), .A2(n2322), .ZN(n2311) );
  NAND2_X1 U1318 ( .A1(NEXT_PC[27]), .A2(n2027), .ZN(n2310) );
  NAND3_X1 U1319 ( .A1(n2312), .A2(n2311), .A3(n2310), .ZN(PRED[27]) );
  NAND2_X1 U1320 ( .A1(PRED_TK[28]), .A2(n1996), .ZN(n2315) );
  NAND2_X1 U1321 ( .A1(NEW_PC[28]), .A2(n2322), .ZN(n2314) );
  NAND2_X1 U1322 ( .A1(NEXT_PC[28]), .A2(n2323), .ZN(n2313) );
  NAND3_X1 U1323 ( .A1(n2315), .A2(n2314), .A3(n2313), .ZN(PRED[28]) );
  NAND2_X1 U1324 ( .A1(PRED_TK[29]), .A2(n1996), .ZN(n2318) );
  NAND2_X1 U1325 ( .A1(NEW_PC[29]), .A2(n2322), .ZN(n2317) );
  NAND2_X1 U1326 ( .A1(NEXT_PC[29]), .A2(n2027), .ZN(n2316) );
  NAND3_X1 U1327 ( .A1(n2318), .A2(n2317), .A3(n2316), .ZN(PRED[29]) );
  NAND2_X1 U1332 ( .A1(NEW_PC[31]), .A2(n2322), .ZN(n2325) );
  NAND2_X1 U1333 ( .A1(NEXT_PC[31]), .A2(n2027), .ZN(n2324) );
  BP_NB32_BP_LEN4_0_DW01_cmp6_0 eq_100 ( .A({\PRED_HISTORY[1][31] , 
        \PRED_HISTORY[1][30] , \PRED_HISTORY[1][29] , \PRED_HISTORY[1][28] , 
        \PRED_HISTORY[1][27] , \PRED_HISTORY[1][26] , \PRED_HISTORY[1][25] , 
        \PRED_HISTORY[1][24] , \PRED_HISTORY[1][23] , \PRED_HISTORY[1][22] , 
        \PRED_HISTORY[1][21] , \PRED_HISTORY[1][20] , \PRED_HISTORY[1][19] , 
        \PRED_HISTORY[1][18] , \PRED_HISTORY[1][17] , \PRED_HISTORY[1][16] , 
        \PRED_HISTORY[1][15] , \PRED_HISTORY[1][14] , \PRED_HISTORY[1][13] , 
        \PRED_HISTORY[1][12] , \PRED_HISTORY[1][11] , \PRED_HISTORY[1][10] , 
        \PRED_HISTORY[1][9] , \PRED_HISTORY[1][8] , \PRED_HISTORY[1][7] , 
        \PRED_HISTORY[1][6] , \PRED_HISTORY[1][5] , \PRED_HISTORY[1][4] , 
        \PRED_HISTORY[1][3] , \PRED_HISTORY[1][2] , \PRED_HISTORY[1][1] , 
        \PRED_HISTORY[1][0] }), .B(EX_PC), .TC(1'b0), .EQ(N815) );
  BP_NB32_BP_LEN4_0_DW01_cmp6_1 eq_59 ( .A({N90, N91, N92, N93, N94, N95, N96, 
        N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, 
        N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, 
        N121}), .B(CURR_PC), .TC(1'b0), .EQ(N122) );
  BP_NB32_BP_LEN4_0_DW01_add_1 add_49_2 ( .A(NEXT_PC), .B({INST[15], INST[15], 
        INST[15], INST[15], INST[15], INST[15], INST[15], INST[15], INST[15], 
        INST[15], INST[15], INST[15], INST[15], INST[15], INST[15], INST[15], 
        INST[15:0]}), .CI(1'b0), .SUM(PRED_TK) );
  DFFR_X2 \PRED_HISTORY_reg[0][23]  ( .D(PRED[23]), .CK(CLK), .RN(n2209), .Q(
        \PRED_HISTORY[0][23] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][30]  ( .D(PRED[30]), .CK(CLK), .RN(n2208), .Q(
        \PRED_HISTORY[0][30] ) );
  NOR2_X1 U1151 ( .A1(n747), .A2(n749), .ZN(n57) );
  CLKBUF_X1 U74 ( .A(N815), .Z(n1963) );
  NOR2_X1 U1334 ( .A1(N815), .A2(n749), .ZN(MISS_HIT[0]) );
  INV_X1 U1198 ( .A(N122), .ZN(n2217) );
  NAND2_X1 U126 ( .A1(n2366), .A2(n2221), .ZN(n2027) );
  INV_X1 U1206 ( .A(n2223), .ZN(n2219) );
  MUX2_X1 U1208 ( .A(n2223), .B(n2222), .S(n2330), .Z(n2221) );
  NAND2_X2 U1202 ( .A1(n2217), .A2(n2330), .ZN(n2366) );
  INV_X1 U1201 ( .A(n2224), .ZN(n2330) );
  BUF_X1 U136 ( .A(n1965), .Z(n1995) );
  NAND2_X1 U73 ( .A1(PRED_TK[31]), .A2(n1965), .ZN(n2326) );
  BUF_X1 U135 ( .A(n1965), .Z(n1994) );
  AND3_X1 U243 ( .A1(N122), .A2(n2330), .A3(n2222), .ZN(n1965) );
  NAND2_X1 U125 ( .A1(n2366), .A2(n2221), .ZN(n2323) );
  OAI221_X1 U1219 ( .B1(n2237), .B2(n2236), .C1(n2235), .C2(n2234), .A(n2233), 
        .ZN(PRED[2]) );
  NOR2_X1 U1088 ( .A1(n2237), .A2(n2229), .ZN(n2230) );
  NOR2_X1 U1087 ( .A1(n2237), .A2(n2225), .ZN(n2226) );
  NAND2_X1 U160 ( .A1(n2224), .A2(n2223), .ZN(n2237) );
  BUF_X1 U138 ( .A(n1965), .Z(n1996) );
  NAND2_X1 U1328 ( .A1(PRED_TK[30]), .A2(n1996), .ZN(n2321) );
  NAND2_X1 U1330 ( .A1(NEXT_PC[30]), .A2(n2323), .ZN(n2319) );
  INV_X4 U65 ( .A(n2237), .ZN(n2322) );
  NAND2_X1 U1329 ( .A1(NEW_PC[30]), .A2(n2322), .ZN(n2320) );
  NAND2_X1 U66 ( .A1(n2321), .A2(n2368), .ZN(PRED[30]) );
  INV_X1 U1331 ( .A(n2367), .ZN(n2368) );
  NAND2_X1 U1338 ( .A1(n2319), .A2(n2320), .ZN(n2367) );
endmodule


module FD_INJ_NB32_4 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n1, n34, n35;
  wire   [31:0] TMP_D;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n35), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n35), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n34), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n34), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n34), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n34), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n1), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n1), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n1), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n1), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n1), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n1), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n1), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n1), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n1), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n1), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n1), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n1), .Q(Q[0]) );
  BUF_X1 U3 ( .A(RESET), .Z(n1) );
  BUF_X1 U4 ( .A(RESET), .Z(n34) );
  BUF_X1 U5 ( .A(RESET), .Z(n35) );
  AND2_X1 U6 ( .A1(D[4]), .A2(INJ_ZERO), .ZN(TMP_D[4]) );
  AND2_X1 U7 ( .A1(D[6]), .A2(INJ_ZERO), .ZN(TMP_D[6]) );
  AND2_X1 U8 ( .A1(D[7]), .A2(INJ_ZERO), .ZN(TMP_D[7]) );
  AND2_X1 U9 ( .A1(D[5]), .A2(INJ_ZERO), .ZN(TMP_D[5]) );
  AND2_X1 U10 ( .A1(D[8]), .A2(INJ_ZERO), .ZN(TMP_D[8]) );
  AND2_X1 U11 ( .A1(D[10]), .A2(INJ_ZERO), .ZN(TMP_D[10]) );
  AND2_X1 U12 ( .A1(D[11]), .A2(INJ_ZERO), .ZN(TMP_D[11]) );
  AND2_X1 U13 ( .A1(D[12]), .A2(INJ_ZERO), .ZN(TMP_D[12]) );
  AND2_X1 U14 ( .A1(D[13]), .A2(INJ_ZERO), .ZN(TMP_D[13]) );
  AND2_X1 U15 ( .A1(D[14]), .A2(INJ_ZERO), .ZN(TMP_D[14]) );
  AND2_X1 U16 ( .A1(D[16]), .A2(INJ_ZERO), .ZN(TMP_D[16]) );
  AND2_X1 U17 ( .A1(D[17]), .A2(INJ_ZERO), .ZN(TMP_D[17]) );
  AND2_X1 U18 ( .A1(D[18]), .A2(INJ_ZERO), .ZN(TMP_D[18]) );
  AND2_X1 U19 ( .A1(D[19]), .A2(INJ_ZERO), .ZN(TMP_D[19]) );
  AND2_X1 U20 ( .A1(D[20]), .A2(INJ_ZERO), .ZN(TMP_D[20]) );
  AND2_X1 U21 ( .A1(D[22]), .A2(INJ_ZERO), .ZN(TMP_D[22]) );
  AND2_X1 U22 ( .A1(D[23]), .A2(INJ_ZERO), .ZN(TMP_D[23]) );
  AND2_X1 U23 ( .A1(D[24]), .A2(INJ_ZERO), .ZN(TMP_D[24]) );
  AND2_X1 U24 ( .A1(D[26]), .A2(INJ_ZERO), .ZN(TMP_D[26]) );
  AND2_X1 U25 ( .A1(D[28]), .A2(INJ_ZERO), .ZN(TMP_D[28]) );
  AND2_X1 U26 ( .A1(D[21]), .A2(INJ_ZERO), .ZN(TMP_D[21]) );
  AND2_X1 U27 ( .A1(D[25]), .A2(INJ_ZERO), .ZN(TMP_D[25]) );
  AND2_X1 U28 ( .A1(D[29]), .A2(INJ_ZERO), .ZN(TMP_D[29]) );
  AND2_X1 U29 ( .A1(D[30]), .A2(INJ_ZERO), .ZN(TMP_D[30]) );
  AND2_X1 U30 ( .A1(D[15]), .A2(INJ_ZERO), .ZN(TMP_D[15]) );
  AND2_X1 U31 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
  AND2_X1 U32 ( .A1(INJ_ZERO), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U33 ( .A1(D[3]), .A2(INJ_ZERO), .ZN(TMP_D[3]) );
  AND2_X1 U34 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U35 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U36 ( .A1(D[31]), .A2(INJ_ZERO), .ZN(TMP_D[31]) );
  AND2_X1 U37 ( .A1(D[27]), .A2(INJ_ZERO), .ZN(TMP_D[27]) );
endmodule


module FD_INJ_NB1_1 ( CK, RESET, INJ_ZERO, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   \TMP_D[0] ;

  DFFR_X1 \Q_reg[0]  ( .D(\TMP_D[0] ), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[0]), .ZN(\TMP_D[0] ) );
endmodule


module FD_INJ_NB1_2 ( CK, RESET, INJ_ZERO, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   \TMP_D[0] ;

  DFFR_X1 \Q_reg[0]  ( .D(\TMP_D[0] ), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[0]), .ZN(\TMP_D[0] ) );
endmodule


module FD_NB2_2 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB4_0 ( CK, RESET, D, Q );
  input [3:0] D;
  output [3:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB3_0 ( CK, RESET, D, Q );
  input [2:0] D;
  output [2:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB4_1 ( CK, RESET, D, Q );
  input [3:0] D;
  output [3:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB3_1 ( CK, RESET, D, Q );
  input [2:0] D;
  output [2:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB2_3 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_21 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_22 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB11_0 ( CK, RESET, D, Q );
  input [10:0] D;
  output [10:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(RESET), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(RESET), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(RESET), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(RESET), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(RESET), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB11_1 ( CK, RESET, D, Q );
  input [10:0] D;
  output [10:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(RESET), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(RESET), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(RESET), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(RESET), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(RESET), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_2 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_3 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FOREWARD_UNIT_NB32_LS5_0 ( .INST_EX({\INST_EX[1] , \INST_EX[0] }), 
    .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }), INST_T_EX, Rs_EX, Rt_EX, Rd_MEM, 
        Rd_WB, CTL_MUX1, CTL_MUX2 );
  input [4:0] Rs_EX;
  input [4:0] Rt_EX;
  input [4:0] Rd_MEM;
  input [4:0] Rd_WB;
  output [1:0] CTL_MUX1;
  output [1:0] CTL_MUX2;
  input \INST_EX[1] , \INST_EX[0] , \INST_MEM[1] , \INST_MEM[0] , INST_T_EX;
  wire   n2, n3, n4, n5, n24, n25, n26, n27, n28, n29, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         net415672, net417563, n8, n7, n40, n39, n38, n37, n36, n35, n34, n33,
         n32, n31, n30, n23, n22, n21, n20, n19, n18, n17, n1, n41, n16, n14,
         n13, net428936, net428935, net428928, n61, n62;
  assign n2 = Rd_MEM[1];

  NAND2_X1 U9 ( .A1(n4), .A2(n5), .ZN(n54) );
  AND4_X2 U10 ( .A1(n59), .A2(n60), .A3(n58), .A4(n57), .ZN(CTL_MUX1[1]) );
  NAND2_X1 U14 ( .A1(n29), .A2(n28), .ZN(n50) );
  NOR2_X1 U35 ( .A1(Rd_WB[0]), .A2(Rd_WB[1]), .ZN(n25) );
  NAND3_X1 U37 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n29) );
  INV_X1 U38 ( .A(INST_MEM[0]), .ZN(n27) );
  NAND2_X1 U39 ( .A1(INST_MEM[1]), .A2(n27), .ZN(n28) );
  XOR2_X1 U46 ( .A(Rs_EX[4]), .B(n3), .Z(n42) );
  NAND2_X1 U52 ( .A1(n43), .A2(n44), .ZN(n45) );
  NOR2_X1 U53 ( .A1(n46), .A2(n45), .ZN(n47) );
  NAND3_X1 U54 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n59) );
  INV_X1 U55 ( .A(n59), .ZN(CTL_MUX1[0]) );
  INV_X1 U56 ( .A(n50), .ZN(n60) );
  XNOR2_X1 U58 ( .A(Rs_EX[3]), .B(Rd_WB[3]), .ZN(n51) );
  AND2_X1 U59 ( .A1(n52), .A2(n51), .ZN(n58) );
  XOR2_X1 U60 ( .A(Rs_EX[0]), .B(Rd_WB[0]), .Z(n56) );
  XNOR2_X1 U61 ( .A(Rs_EX[1]), .B(Rd_WB[1]), .ZN(n53) );
  NAND2_X1 U62 ( .A1(n54), .A2(n53), .ZN(n55) );
  NOR2_X1 U63 ( .A1(n56), .A2(n55), .ZN(n57) );
  OR2_X1 U6 ( .A1(Rs_EX[2]), .A2(Rd_WB[2]), .ZN(n5) );
  NAND2_X1 U8 ( .A1(Rs_EX[2]), .A2(Rd_WB[2]), .ZN(n4) );
  INV_X1 U34 ( .A(Rd_WB[2]), .ZN(n26) );
  XNOR2_X1 U57 ( .A(Rd_WB[4]), .B(Rs_EX[4]), .ZN(n52) );
  NOR2_X1 U36 ( .A1(Rd_WB[3]), .A2(Rd_WB[4]), .ZN(n24) );
  NAND2_X1 U29 ( .A1(n18), .A2(n17), .ZN(n19) );
  NOR2_X1 U30 ( .A1(n19), .A2(n20), .ZN(n21) );
  XNOR2_X1 U48 ( .A(n1), .B(Rs_EX[3]), .ZN(n48) );
  XNOR2_X1 U25 ( .A(Rt_EX[3]), .B(n1), .ZN(n22) );
  NAND3_X1 U31 ( .A1(n23), .A2(n21), .A3(n22), .ZN(n40) );
  NOR2_X1 U16 ( .A1(n30), .A2(n40), .ZN(CTL_MUX2[0]) );
  INV_X1 U32 ( .A(INST_T_EX), .ZN(n30) );
  NOR2_X1 U15 ( .A1(n50), .A2(n30), .ZN(n38) );
  XNOR2_X1 U40 ( .A(Rd_WB[1]), .B(Rt_EX[1]), .ZN(n32) );
  XNOR2_X1 U41 ( .A(Rd_WB[0]), .B(Rt_EX[0]), .ZN(n31) );
  NAND2_X1 U42 ( .A1(n32), .A2(n31), .ZN(n36) );
  OR2_X1 U7 ( .A1(Rd_WB[3]), .A2(Rt_EX[3]), .ZN(n8) );
  NAND2_X1 U11 ( .A1(Rd_WB[3]), .A2(Rt_EX[3]), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n8), .A2(n7), .ZN(n34) );
  XNOR2_X1 U43 ( .A(Rd_WB[2]), .B(Rt_EX[2]), .ZN(n33) );
  NAND2_X1 U44 ( .A1(n33), .A2(n34), .ZN(n35) );
  NOR2_X1 U45 ( .A1(n36), .A2(n35), .ZN(n37) );
  XNOR2_X1 U33 ( .A(Rd_WB[4]), .B(Rt_EX[4]), .ZN(n39) );
  AND4_X2 U5 ( .A1(n40), .A2(n38), .A3(n37), .A4(n39), .ZN(CTL_MUX2[1]) );
  INV_X1 U22 ( .A(INST_EX[0]), .ZN(n13) );
  NAND2_X1 U23 ( .A1(n13), .A2(INST_EX[1]), .ZN(n14) );
  NOR2_X1 U24 ( .A1(n41), .A2(n16), .ZN(n23) );
  NOR2_X1 U47 ( .A1(n42), .A2(n41), .ZN(n49) );
  NAND3_X1 syn154 ( .A1(n62), .A2(net428936), .A3(net428935), .ZN(net428928)
         );
  BUF_X1 U2 ( .A(Rd_MEM[2]), .Z(n61) );
  NAND2_X1 U3 ( .A1(net428928), .A2(n14), .ZN(n41) );
  NOR2_X1 U4 ( .A1(Rd_MEM[4]), .A2(Rd_MEM[3]), .ZN(net428935) );
  INV_X1 U13 ( .A(Rd_MEM[2]), .ZN(net428936) );
  NOR2_X1 U17 ( .A1(Rd_MEM[0]), .A2(n2), .ZN(n62) );
  XOR2_X1 U18 ( .A(Rd_MEM[4]), .B(Rt_EX[4]), .Z(n16) );
  CLKBUF_X1 U19 ( .A(Rd_MEM[4]), .Z(n3) );
  CLKBUF_X1 U20 ( .A(Rd_MEM[3]), .Z(n1) );
  XNOR2_X1 U21 ( .A(Rd_MEM[2]), .B(Rt_EX[2]), .ZN(n18) );
  XNOR2_X1 U26 ( .A(n61), .B(Rs_EX[2]), .ZN(n44) );
  XNOR2_X1 U27 ( .A(n2), .B(Rt_EX[1]), .ZN(n17) );
  CLKBUF_X1 U28 ( .A(n2), .Z(net417563) );
  XOR2_X1 U49 ( .A(Rd_MEM[0]), .B(Rt_EX[0]), .Z(n20) );
  CLKBUF_X1 U50 ( .A(Rd_MEM[0]), .Z(net415672) );
  XNOR2_X1 U51 ( .A(net417563), .B(Rs_EX[1]), .ZN(n43) );
  XOR2_X1 U64 ( .A(Rs_EX[0]), .B(net415672), .Z(n46) );
endmodule


module WRITE_BACK_UNIT_NB32_LS5_0 ( MEM_ALU_SEL, DEST_IN, FROM_ALU, FROM_MEM, 
        DATA_OUT, DEST_OUT );
  input [4:0] DEST_IN;
  input [31:0] FROM_ALU;
  input [31:0] FROM_MEM;
  output [31:0] DATA_OUT;
  output [4:0] DEST_OUT;
  input MEM_ALU_SEL;

  assign DEST_OUT[4] = DEST_IN[4];
  assign DEST_OUT[3] = DEST_IN[3];
  assign DEST_OUT[2] = DEST_IN[2];
  assign DEST_OUT[1] = DEST_IN[1];
  assign DEST_OUT[0] = DEST_IN[0];

  MUX21_generic_NB32_0 wb_mux ( .A(FROM_ALU), .B(FROM_MEM), .SEL(MEM_ALU_SEL), 
        .Y(DATA_OUT) );
endmodule


module MEMORY_UNIT_NB32_LS5_0 ( CLK, RST, DEST_IN, FROM_MEM, FROM_ALU, ALU_OUT, 
        MEM_OUT, DEST_OUT );
  input [4:0] DEST_IN;
  input [31:0] FROM_MEM;
  input [31:0] FROM_ALU;
  output [31:0] ALU_OUT;
  output [31:0] MEM_OUT;
  output [4:0] DEST_OUT;
  input CLK, RST;


  FD_NB32_1 exec_reg ( .CK(CLK), .RESET(RST), .D(FROM_ALU), .Q(ALU_OUT) );
  FD_NB32_0 mem_reg ( .CK(CLK), .RESET(RST), .D(FROM_MEM), .Q(MEM_OUT) );
  FD_NB5_0 dest_reg ( .CK(CLK), .RESET(RST), .D(DEST_IN), .Q(DEST_OUT) );
endmodule


module EXECUTION_UNIT_NB32_LS5_0 ( FW_MUX1_SEL, FW_MUX2_SEL, FW_EX, FW_MEM, A, 
        B, C, D, DEST_IN, CLK, RST, US, MUX1_SEL, MUX2_SEL, UN_SEL, OP_SEL, 
        US_MEM, TEMP_PC, ALU_OUT, IMM_OUT, DEST_OUT );
  input [1:0] FW_MUX1_SEL;
  input [1:0] FW_MUX2_SEL;
  input [31:0] FW_EX;
  input [31:0] FW_MEM;
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [4:0] DEST_IN;
  input [2:0] UN_SEL;
  input [3:0] OP_SEL;
  output [31:0] TEMP_PC;
  output [31:0] ALU_OUT;
  output [31:0] IMM_OUT;
  output [4:0] DEST_OUT;
  input CLK, RST, US, MUX1_SEL, MUX2_SEL;
  output US_MEM;
  wire   CA_OUT, n7, n8, n1, n2, n3, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;
  wire   [30:0] TERM1;
  wire   [30:0] TERM2;
  wire   [1:0] MSB;
  wire   [31:0] TERM4;
  wire   [31:0] TERM5;
  wire   [31:0] TERM3;
  wire   [31:0] MUL_OUT;
  wire   [31:0] SHFT_OUT;
  wire   [31:0] COMP_OUT;
  wire   [31:0] LOGIC_OUT;
  wire   [4:0] TMP_DEST_OUT;
  wire   [31:0] MUX2_OUT;
  wire   [31:0] JMP_RET;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  BUF_X2 U4 ( .A(TERM1[13]), .Z(n35) );
  CLKBUF_X1 U7 ( .A(TERM2[8]), .Z(n1) );
  CLKBUF_X1 U8 ( .A(TEMP_PC[20]), .Z(n2) );
  BUF_X2 U9 ( .A(TERM1[9]), .Z(n31) );
  XNOR2_X1 U10 ( .A(TERM2[4]), .B(n41), .ZN(TERM3[4]) );
  CLKBUF_X1 U11 ( .A(TERM2[5]), .Z(n15) );
  CLKBUF_X1 U12 ( .A(TERM2[7]), .Z(n3) );
  CLKBUF_X1 U13 ( .A(TERM2[2]), .Z(n9) );
  CLKBUF_X1 U14 ( .A(TERM2[14]), .Z(n10) );
  CLKBUF_X1 U15 ( .A(TERM2[10]), .Z(n11) );
  CLKBUF_X1 U16 ( .A(TERM1[6]), .Z(n29) );
  BUF_X4 U17 ( .A(TERM1[10]), .Z(n32) );
  CLKBUF_X1 U18 ( .A(TERM1[15]), .Z(n36) );
  CLKBUF_X1 U19 ( .A(TERM1[11]), .Z(n33) );
  CLKBUF_X1 U20 ( .A(TERM2[6]), .Z(n12) );
  CLKBUF_X1 U21 ( .A(TEMP_PC[27]), .Z(n13) );
  CLKBUF_X1 U22 ( .A(TERM1[5]), .Z(n28) );
  CLKBUF_X1 U23 ( .A(TERM2[3]), .Z(n14) );
  CLKBUF_X1 U24 ( .A(TERM2[15]), .Z(n16) );
  CLKBUF_X1 U25 ( .A(TEMP_PC[21]), .Z(n17) );
  BUF_X1 U26 ( .A(TERM2[12]), .Z(n18) );
  CLKBUF_X1 U27 ( .A(TEMP_PC[29]), .Z(n19) );
  XNOR2_X1 U28 ( .A(TERM2[5]), .B(n41), .ZN(TERM3[5]) );
  CLKBUF_X3 U30 ( .A(TERM1[12]), .Z(n34) );
  CLKBUF_X3 U31 ( .A(TERM1[8]), .Z(n30) );
  AND3_X1 U32 ( .A1(OP_SEL[2]), .A2(n38), .A3(n8), .ZN(n7) );
  NOR2_X1 U33 ( .A1(OP_SEL[3]), .A2(OP_SEL[1]), .ZN(n8) );
  OR2_X1 U34 ( .A1(n7), .A2(DEST_IN[0]), .ZN(TMP_DEST_OUT[0]) );
  OR2_X1 U35 ( .A1(n7), .A2(DEST_IN[1]), .ZN(TMP_DEST_OUT[1]) );
  OR2_X1 U36 ( .A1(n7), .A2(DEST_IN[2]), .ZN(TMP_DEST_OUT[2]) );
  OR2_X1 U37 ( .A1(n7), .A2(DEST_IN[3]), .ZN(TMP_DEST_OUT[3]) );
  OR2_X1 U38 ( .A1(n7), .A2(DEST_IN[4]), .ZN(TMP_DEST_OUT[4]) );
  NAND2_X1 U40 ( .A1(TERM2[3]), .A2(n41), .ZN(n22) );
  NAND2_X1 U41 ( .A1(n20), .A2(n21), .ZN(n23) );
  NAND2_X1 U42 ( .A1(n23), .A2(n22), .ZN(TERM3[3]) );
  INV_X1 U43 ( .A(TERM2[3]), .ZN(n20) );
  INV_X1 U44 ( .A(n41), .ZN(n21) );
  BUF_X2 U46 ( .A(TERM1[1]), .Z(n27) );
  XNOR2_X1 U47 ( .A(TERM2[6]), .B(n41), .ZN(TERM3[6]) );
  XNOR2_X1 U48 ( .A(TERM2[13]), .B(n40), .ZN(TERM3[13]) );
  XNOR2_X1 U50 ( .A(TERM2[9]), .B(n40), .ZN(TERM3[9]) );
  XNOR2_X1 U51 ( .A(TERM2[2]), .B(n41), .ZN(TERM3[2]) );
  XNOR2_X1 U52 ( .A(TERM2[1]), .B(n41), .ZN(TERM3[1]) );
  CLKBUF_X1 U53 ( .A(TERM1[0]), .Z(n26) );
  CLKBUF_X1 U54 ( .A(TEMP_PC[25]), .Z(n25) );
  INV_X2 U55 ( .A(n38), .ZN(n39) );
  INV_X2 U56 ( .A(n38), .ZN(n40) );
  XNOR2_X1 U58 ( .A(MSB[0]), .B(n39), .ZN(TERM3[31]) );
  XNOR2_X1 U59 ( .A(TERM2[30]), .B(n39), .ZN(TERM3[30]) );
  XNOR2_X1 U60 ( .A(TERM2[29]), .B(n39), .ZN(TERM3[29]) );
  XNOR2_X1 U61 ( .A(TERM2[28]), .B(n39), .ZN(TERM3[28]) );
  XNOR2_X1 U62 ( .A(TERM2[27]), .B(n39), .ZN(TERM3[27]) );
  XNOR2_X1 U63 ( .A(TERM2[26]), .B(n39), .ZN(TERM3[26]) );
  XNOR2_X1 U64 ( .A(TERM2[25]), .B(n39), .ZN(TERM3[25]) );
  XNOR2_X1 U65 ( .A(TERM2[24]), .B(n39), .ZN(TERM3[24]) );
  XNOR2_X1 U66 ( .A(TERM2[23]), .B(n39), .ZN(TERM3[23]) );
  XNOR2_X1 U67 ( .A(TERM2[22]), .B(n39), .ZN(TERM3[22]) );
  XNOR2_X1 U68 ( .A(TERM2[21]), .B(n39), .ZN(TERM3[21]) );
  XNOR2_X1 U69 ( .A(TERM2[20]), .B(n39), .ZN(TERM3[20]) );
  XNOR2_X1 U70 ( .A(TERM2[19]), .B(n40), .ZN(TERM3[19]) );
  XNOR2_X1 U71 ( .A(TERM2[18]), .B(n40), .ZN(TERM3[18]) );
  XNOR2_X1 U72 ( .A(TERM2[17]), .B(n40), .ZN(TERM3[17]) );
  XNOR2_X1 U73 ( .A(TERM2[16]), .B(n40), .ZN(TERM3[16]) );
  XNOR2_X1 U74 ( .A(TERM2[15]), .B(n40), .ZN(TERM3[15]) );
  XNOR2_X1 U75 ( .A(TERM2[14]), .B(n40), .ZN(TERM3[14]) );
  XNOR2_X1 U76 ( .A(TERM2[12]), .B(n40), .ZN(TERM3[12]) );
  XNOR2_X1 U77 ( .A(TERM2[11]), .B(n40), .ZN(TERM3[11]) );
  XNOR2_X1 U78 ( .A(TERM2[10]), .B(n40), .ZN(TERM3[10]) );
  XNOR2_X1 U79 ( .A(TERM2[8]), .B(n40), .ZN(TERM3[8]) );
  XNOR2_X1 U80 ( .A(TERM2[7]), .B(n41), .ZN(TERM3[7]) );
  MUX21_generic_NB32_2 mux1 ( .A(A), .B(D), .SEL(MUX1_SEL), .Y(TERM4) );
  MUX21_generic_NB32_1 mux2 ( .A(B), .B(C), .SEL(MUX2_SEL), .Y(TERM5) );
  MUX31_generic_NB32_1 fW_mux1 ( .A(TERM4), .B(FW_EX), .C(FW_MEM), .SEL(
        FW_MUX1_SEL), .Y({MSB[1], TERM1}) );
  MUX31_generic_NB32_0 fw_mux2 ( .A(TERM5), .B(FW_EX), .C(FW_MEM), .SEL(
        FW_MUX2_SEL), .Y({MSB[0], TERM2}) );
  p4addgen_NB32_CW4_8 adder ( .A({MSB[1], TERM1[30:14], n35, n34, TERM1[11], 
        n32, n31, n30, TERM1[7:2], n27, TERM1[0]}), .B(TERM3), .Ci(n38), .Co(
        CA_OUT), .S(TEMP_PC) );
  BOOTHMUL_NB32_0 multiplier ( .A({n36, TERM1[14], n35, n34, n33, n32, n31, 
        n30, TERM1[7], n29, n28, TERM1[4:2], n27, n26}), .B({n16, n10, n42, 
        n18, n43, n11, TERM2[9], n1, n3, n12, n15, TERM2[4], n14, n9, TERM2[1], 
        n24}), .C(MUL_OUT) );
  SHIFTER_NB32_LS5_0 shift_rot ( .FUNC({OP_SEL[1], n37}), .US(US), .DATA1({
        MSB[1], TERM1[30:14], n35, n34, n33, n32, n31, n30, TERM1[7], n29, n28, 
        TERM1[4:2], n27, n26}), .DATA2({TERM2[4], n14, n9, TERM2[1], n24}), 
        .OUTSHFT(SHFT_OUT) );
  COMPARATOR_NB32_0 comparison ( .AdderRes({TEMP_PC[31:30], n19, TEMP_PC[28], 
        n13, n45, n25, TEMP_PC[24:22], n17, n2, TEMP_PC[19:15], n44, 
        TEMP_PC[13:0]}), .MSB(MSB), .CO(CA_OUT), .OP_CODE(OP_SEL[3:1]), .US(US), .SOUT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, COMP_OUT[0]}) );
  LOGIC_NB32_0 log_un ( .SEL({OP_SEL[3:1], n37}), .A({MSB[1], TERM1[30:16], 
        n36, TERM1[14], n35, n34, n33, n32, n31, n30, TERM1[7], n29, n28, 
        TERM1[4:2], n27, n26}), .B({MSB[0], TERM2[30:15], n10, TERM2[13], n18, 
        TERM2[11], n11, TERM2[9], n1, n3, n12, n15, TERM2[4], n14, n9, 
        TERM2[1], n24}), .RES(LOGIC_OUT) );
  FD_NB5_1 destination_register ( .CK(CLK), .RESET(RST), .D(TMP_DEST_OUT), .Q(
        DEST_OUT) );
  FD_NB32_3 output_register ( .CK(CLK), .RESET(RST), .D(MUX2_OUT), .Q(ALU_OUT)
         );
  FD_NB32_2 imm_register ( .CK(CLK), .RESET(RST), .D(B), .Q(IMM_OUT) );
  FD_NB1_0 us_register ( .CK(CLK), .RESET(RST), .D(US), .Q(US_MEM) );
  MUX61_generic_NB32_0 mux_out ( .A({TEMP_PC[31:30], n19, TEMP_PC[28], n13, 
        n45, n25, TEMP_PC[24:22], n17, n2, TEMP_PC[19:0]}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, COMP_OUT[0]}), .C(MUL_OUT), .D(SHFT_OUT), 
        .E(LOGIC_OUT), .F(JMP_RET), .SEL(UN_SEL), .Y(MUX2_OUT) );
  EXECUTION_UNIT_NB32_LS5_0_DW01_add_0 add_202 ( .A(D), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(JMP_RET) );
  CLKBUF_X1 U39 ( .A(OP_SEL[0]), .Z(n37) );
  CLKBUF_X1 U49 ( .A(TERM2[0]), .Z(n24) );
  CLKBUF_X2 U57 ( .A(OP_SEL[0]), .Z(n38) );
  INV_X2 U45 ( .A(n38), .ZN(n41) );
  XNOR2_X1 U29 ( .A(TERM2[0]), .B(n41), .ZN(TERM3[0]) );
  CLKBUF_X1 U112 ( .A(TERM2[13]), .Z(n42) );
  CLKBUF_X1 U113 ( .A(TERM2[11]), .Z(n43) );
  CLKBUF_X1 U114 ( .A(TEMP_PC[14]), .Z(n44) );
  CLKBUF_X1 U115 ( .A(TEMP_PC[26]), .Z(n45) );
endmodule


module DECODE_UNIT_NB32_LS5_0 ( CLK, RST, FLUSH, DATAIN, IMM1, IMM2, BR_TYPE, 
        JMP, RI, US, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DEST_IN, HAZARD, 
        US_TO_EX, A, B, C, D, RT, RS, DEST_OUT );
  input [31:0] DATAIN;
  input [25:0] IMM1;
  input [31:0] IMM2;
  input [1:0] BR_TYPE;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [4:0] DEST_IN;
  output [31:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [4:0] RT;
  output [4:0] RS;
  output [4:0] DEST_OUT;
  input CLK, RST, FLUSH, JMP, RI, US, RD1, RD2, WR;
  output HAZARD, US_TO_EX;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n1, n15, n16,
         n17;
  wire   [31:0] OUT1;
  wire   [31:0] OUT2;
  wire   [31:0] EXT1;
  wire   [31:0] TO_IMM1;
  wire   [4:0] DEST_ADD;

  BUF_X2 U2 ( .A(RST), .Z(n17) );
  NOR4_X1 U3 ( .A1(OUT1[23]), .A2(OUT1[22]), .A3(OUT1[21]), .A4(OUT1[20]), 
        .ZN(n10) );
  NOR4_X1 U4 ( .A1(OUT1[9]), .A2(OUT1[8]), .A3(OUT1[7]), .A4(OUT1[6]), .ZN(n14) );
  NOR4_X1 U5 ( .A1(OUT1[5]), .A2(OUT1[4]), .A3(OUT1[3]), .A4(OUT1[31]), .ZN(
        n13) );
  NOR4_X1 U6 ( .A1(OUT1[30]), .A2(OUT1[2]), .A3(OUT1[29]), .A4(OUT1[28]), .ZN(
        n12) );
  NOR4_X1 U7 ( .A1(OUT1[27]), .A2(OUT1[26]), .A3(OUT1[25]), .A4(OUT1[24]), 
        .ZN(n11) );
  NAND4_X1 U8 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n6) );
  NOR4_X1 U9 ( .A1(OUT1[12]), .A2(OUT1[11]), .A3(OUT1[10]), .A4(OUT1[0]), .ZN(
        n7) );
  NOR4_X1 U10 ( .A1(OUT1[16]), .A2(OUT1[15]), .A3(OUT1[14]), .A4(OUT1[13]), 
        .ZN(n8) );
  NOR4_X1 U11 ( .A1(OUT1[1]), .A2(OUT1[19]), .A3(OUT1[18]), .A4(OUT1[17]), 
        .ZN(n9) );
  AND2_X1 U12 ( .A1(EXT1[25]), .A2(n15), .ZN(TO_IMM1[25]) );
  AND2_X1 U13 ( .A1(EXT1[26]), .A2(n15), .ZN(TO_IMM1[26]) );
  AND2_X1 U14 ( .A1(EXT1[27]), .A2(n15), .ZN(TO_IMM1[27]) );
  AND2_X1 U15 ( .A1(EXT1[28]), .A2(n1), .ZN(TO_IMM1[28]) );
  AND2_X1 U16 ( .A1(EXT1[29]), .A2(n1), .ZN(TO_IMM1[29]) );
  AND2_X1 U17 ( .A1(EXT1[30]), .A2(n1), .ZN(TO_IMM1[30]) );
  AND2_X1 U18 ( .A1(EXT1[31]), .A2(n1), .ZN(TO_IMM1[31]) );
  BUF_X1 U19 ( .A(n2), .Z(n15) );
  BUF_X1 U20 ( .A(n2), .Z(n1) );
  BUF_X1 U21 ( .A(n2), .Z(n16) );
  AND2_X1 U22 ( .A1(EXT1[0]), .A2(n16), .ZN(TO_IMM1[0]) );
  AND2_X1 U23 ( .A1(EXT1[1]), .A2(n15), .ZN(TO_IMM1[1]) );
  AND2_X1 U24 ( .A1(EXT1[2]), .A2(n1), .ZN(TO_IMM1[2]) );
  AND2_X1 U25 ( .A1(EXT1[10]), .A2(n16), .ZN(TO_IMM1[10]) );
  AND2_X1 U26 ( .A1(EXT1[11]), .A2(n16), .ZN(TO_IMM1[11]) );
  AND2_X1 U27 ( .A1(EXT1[12]), .A2(n16), .ZN(TO_IMM1[12]) );
  AND2_X1 U28 ( .A1(EXT1[13]), .A2(n16), .ZN(TO_IMM1[13]) );
  AND2_X1 U29 ( .A1(EXT1[14]), .A2(n16), .ZN(TO_IMM1[14]) );
  AND2_X1 U30 ( .A1(EXT1[15]), .A2(n16), .ZN(TO_IMM1[15]) );
  AND2_X1 U31 ( .A1(EXT1[16]), .A2(n16), .ZN(TO_IMM1[16]) );
  AND2_X1 U32 ( .A1(EXT1[17]), .A2(n15), .ZN(TO_IMM1[17]) );
  AND2_X1 U33 ( .A1(EXT1[18]), .A2(n15), .ZN(TO_IMM1[18]) );
  AND2_X1 U34 ( .A1(EXT1[19]), .A2(n15), .ZN(TO_IMM1[19]) );
  AND2_X1 U35 ( .A1(EXT1[20]), .A2(n15), .ZN(TO_IMM1[20]) );
  AND2_X1 U36 ( .A1(EXT1[21]), .A2(n15), .ZN(TO_IMM1[21]) );
  AND2_X1 U37 ( .A1(EXT1[22]), .A2(n15), .ZN(TO_IMM1[22]) );
  AND2_X1 U38 ( .A1(EXT1[23]), .A2(n15), .ZN(TO_IMM1[23]) );
  AND2_X1 U39 ( .A1(EXT1[24]), .A2(n15), .ZN(TO_IMM1[24]) );
  AND2_X1 U40 ( .A1(EXT1[9]), .A2(n1), .ZN(TO_IMM1[9]) );
  AND2_X1 U41 ( .A1(EXT1[3]), .A2(n1), .ZN(TO_IMM1[3]) );
  AND2_X1 U42 ( .A1(EXT1[4]), .A2(n1), .ZN(TO_IMM1[4]) );
  AND2_X1 U43 ( .A1(EXT1[5]), .A2(n1), .ZN(TO_IMM1[5]) );
  AND2_X1 U44 ( .A1(EXT1[6]), .A2(n1), .ZN(TO_IMM1[6]) );
  AND2_X1 U45 ( .A1(EXT1[7]), .A2(n1), .ZN(TO_IMM1[7]) );
  AND2_X1 U46 ( .A1(EXT1[8]), .A2(n1), .ZN(TO_IMM1[8]) );
  NAND2_X1 U47 ( .A1(n3), .A2(BR_TYPE[1]), .ZN(n2) );
  XNOR2_X1 U48 ( .A(BR_TYPE[0]), .B(n4), .ZN(n3) );
  NOR2_X1 U49 ( .A1(n5), .A2(n6), .ZN(n4) );
  NAND4_X1 U50 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .ZN(n5) );
  register_file_NB32_RS32_0 reg_file ( .CLK(CLK), .RESET(n17), .RD1(RD1), 
        .RD2(RD2), .WR(WR), .ADD_WR(ADD_WR), .ADD_RD1(ADD_RD1), .ADD_RD2(
        ADD_RD2), .DATAIN(DATAIN), .HAZARD(HAZARD), .OUT1(OUT1), .OUT2(OUT2)
         );
  FD_INJ_NB32_3 reg_a ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(OUT1), .Q(
        A) );
  FD_INJ_NB32_2 reg_b ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(OUT2), .Q(
        B) );
  SIGN_EXT_NB32_0 exted ( .A(IMM1), .US(US), .JMP(JMP), .Y(EXT1) );
  FD_INJ_NB1_0 us_register ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(US), 
        .Q(US_TO_EX) );
  FD_INJ_NB32_1 imm_reg1 ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(TO_IMM1), .Q(C) );
  FD_INJ_NB32_0 imm_reg2 ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(IMM2), 
        .Q(D) );
  MUX21_generic_NB5_0 mux_dest ( .A(ADD_RD2), .B(DEST_IN), .SEL(RI), .Y(
        DEST_ADD) );
  FD_INJ_NB5_2 dest_reg ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(DEST_ADD), .Q(DEST_OUT) );
  FD_INJ_NB5_1 rs_reg ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(ADD_RD1), 
        .Q(RS) );
  FD_INJ_NB5_0 rt_reg ( .CK(CLK), .RESET(n17), .INJ_ZERO(FLUSH), .D(ADD_RD2), 
        .Q(RT) );
endmodule


module FETCH_UNIT_NB32_LS5_0 ( CLK, STALL, RST, RST_DEC, PC_SEL, JB_INST, 
        IRAM_OUT, FUNC, OPCODE, CURR_PC, NPC, INST_OUT, MISS_HIT );
  input [31:0] JB_INST;
  input [31:0] IRAM_OUT;
  output [10:0] FUNC;
  output [5:0] OPCODE;
  output [31:0] CURR_PC;
  output [31:0] NPC;
  output [31:0] INST_OUT;
  output [1:0] MISS_HIT;
  input CLK, STALL, RST, RST_DEC, PC_SEL;
  wire   \IRAM_OUT[10] , \IRAM_OUT[9] , \IRAM_OUT[8] , \IRAM_OUT[7] ,
         \IRAM_OUT[6] , \IRAM_OUT[5] , \IRAM_OUT[4] , \IRAM_OUT[3] ,
         \IRAM_OUT[2] , \IRAM_OUT[1] , \IRAM_OUT[0] , \IRAM_OUT[31] ,
         \IRAM_OUT[30] , \IRAM_OUT[29] , \IRAM_OUT[28] , \IRAM_OUT[27] ,
         \IRAM_OUT[26] , n20, n21, TMP_RST, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n15, n16, n17, n18, n22, n23, n24, n25, n26;
  wire   [31:0] NEXT_PC;
  wire   [31:0] NEW_PC;
  wire   [31:0] TMP_INST_OUT;
  wire   [31:0] PRED;
  assign FUNC[10] = \IRAM_OUT[10] ;
  assign \IRAM_OUT[10]  = IRAM_OUT[10];
  assign FUNC[9] = \IRAM_OUT[9] ;
  assign \IRAM_OUT[9]  = IRAM_OUT[9];
  assign FUNC[8] = \IRAM_OUT[8] ;
  assign \IRAM_OUT[8]  = IRAM_OUT[8];
  assign FUNC[7] = \IRAM_OUT[7] ;
  assign \IRAM_OUT[7]  = IRAM_OUT[7];
  assign FUNC[6] = \IRAM_OUT[6] ;
  assign \IRAM_OUT[6]  = IRAM_OUT[6];
  assign FUNC[5] = \IRAM_OUT[5] ;
  assign \IRAM_OUT[5]  = IRAM_OUT[5];
  assign FUNC[4] = \IRAM_OUT[4] ;
  assign \IRAM_OUT[4]  = IRAM_OUT[4];
  assign FUNC[3] = \IRAM_OUT[3] ;
  assign \IRAM_OUT[3]  = IRAM_OUT[3];
  assign FUNC[2] = \IRAM_OUT[2] ;
  assign \IRAM_OUT[2]  = IRAM_OUT[2];
  assign FUNC[1] = \IRAM_OUT[1] ;
  assign \IRAM_OUT[1]  = IRAM_OUT[1];
  assign FUNC[0] = \IRAM_OUT[0] ;
  assign \IRAM_OUT[0]  = IRAM_OUT[0];
  assign OPCODE[5] = \IRAM_OUT[31] ;
  assign \IRAM_OUT[31]  = IRAM_OUT[31];
  assign OPCODE[4] = \IRAM_OUT[30] ;
  assign \IRAM_OUT[30]  = IRAM_OUT[30];
  assign OPCODE[3] = \IRAM_OUT[29] ;
  assign \IRAM_OUT[29]  = IRAM_OUT[29];
  assign OPCODE[2] = \IRAM_OUT[28] ;
  assign \IRAM_OUT[28]  = IRAM_OUT[28];
  assign OPCODE[1] = \IRAM_OUT[27] ;
  assign \IRAM_OUT[27]  = IRAM_OUT[27];
  assign OPCODE[0] = \IRAM_OUT[26] ;
  assign \IRAM_OUT[26]  = IRAM_OUT[26];

  DFF_X1 TMP_RST_reg ( .D(RST), .CK(CLK), .Q(TMP_RST) );
  CLKBUF_X1 U3 ( .A(TMP_INST_OUT[8]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(TMP_INST_OUT[12]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(TMP_INST_OUT[13]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(TMP_INST_OUT[3]), .Z(n6) );
  CLKBUF_X1 U8 ( .A(TMP_INST_OUT[9]), .Z(n7) );
  CLKBUF_X1 U9 ( .A(TMP_INST_OUT[11]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(TMP_INST_OUT[14]), .Z(n9) );
  CLKBUF_X1 U11 ( .A(TMP_INST_OUT[0]), .Z(n10) );
  CLKBUF_X1 U12 ( .A(TMP_INST_OUT[1]), .Z(n11) );
  CLKBUF_X1 U13 ( .A(JB_INST[21]), .Z(n12) );
  CLKBUF_X1 U14 ( .A(TMP_INST_OUT[15]), .Z(n13) );
  CLKBUF_X1 U16 ( .A(n20), .Z(CURR_PC[1]) );
  CLKBUF_X1 U17 ( .A(JB_INST[25]), .Z(n15) );
  FD_INJ_NB32_4 N_PC ( .CK(CLK), .RESET(RST), .INJ_ZERO(n16), .D(NEXT_PC), .Q(
        NPC) );
  BP_NB32_BP_LEN4_0 BP_UNIT ( .CLK(CLK), .RST(RST), .EX_PC(JB_INST), .CURR_PC(
        CURR_PC), .NEXT_PC(NEXT_PC), .NEW_PC(NEW_PC), .INST(TMP_INST_OUT), 
        .MISS_HIT({MISS_HIT[1], n21}), .PRED(PRED) );
  FD_NB32_5 PC ( .CK(CLK), .RESET(TMP_RST), .D(PRED), .Q({CURR_PC[31:2], n20, 
        CURR_PC[0]}) );
  MUX21_generic_NB32_4 flush_mux ( .A({\IRAM_OUT[31] , \IRAM_OUT[30] , 
        \IRAM_OUT[29] , \IRAM_OUT[28] , \IRAM_OUT[27] , \IRAM_OUT[26] , 
        IRAM_OUT[25:11], \IRAM_OUT[10] , \IRAM_OUT[9] , \IRAM_OUT[8] , 
        \IRAM_OUT[7] , \IRAM_OUT[6] , \IRAM_OUT[5] , \IRAM_OUT[4] , 
        \IRAM_OUT[3] , \IRAM_OUT[2] , \IRAM_OUT[1] , \IRAM_OUT[0] }), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n17), .Y(TMP_INST_OUT) );
  FD_NB32_4 INST ( .CK(CLK), .RESET(RST), .D({TMP_INST_OUT[31:16], n13, n9, n5, 
        n4, n8, n24, n7, n2, n23, TMP_INST_OUT[6], n26, n25, n6, 
        TMP_INST_OUT[2], n11, n10}), .Q(INST_OUT) );
  MUX21_generic_NB32_3 pc_mux ( .A({JB_INST[31:27], n22, n15, JB_INST[24:22], 
        n12, JB_INST[20:0]}), .B(NEXT_PC), .SEL(PC_SEL), .Y(NEW_PC) );
  FETCH_UNIT_NB32_LS5_0_DW01_add_0 add_123 ( .A({CURR_PC[31:2], n20, 
        CURR_PC[0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), 
        .CI(1'b0), .SUM(NEXT_PC) );
  CLKBUF_X1 U20 ( .A(n21), .Z(MISS_HIT[0]) );
  INV_X1 U15 ( .A(STALL), .ZN(n18) );
  CLKBUF_X1 U18 ( .A(n17), .Z(n16) );
  AOI21_X2 U19 ( .B1(n21), .B2(MISS_HIT[1]), .A(n18), .ZN(n17) );
  CLKBUF_X1 U21 ( .A(JB_INST[26]), .Z(n22) );
  CLKBUF_X1 U22 ( .A(TMP_INST_OUT[7]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(TMP_INST_OUT[10]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(TMP_INST_OUT[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(TMP_INST_OUT[5]), .Z(n26) );
endmodule


module DLX_CU_0 ( CLK, RST, OPCODE, FUNC, FLUSH, STALL, JMP, RI, BR_TYPE, RD1, 
        RD2, US, MUX1_SEL, MUX2_SEL, UN_SEL, OP_SEL, PC_SEL, RW, D_TYPE, WR, 
        MEM_ALU_SEL, INST_T_EX, .INST_EX({\INST_EX[1] , \INST_EX[0] }), 
    .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }) );
  input [5:0] OPCODE;
  input [10:0] FUNC;
  output [1:0] BR_TYPE;
  output [2:0] UN_SEL;
  output [3:0] OP_SEL;
  output [1:0] D_TYPE;
  input CLK, RST, FLUSH;
  output STALL, JMP, RI, RD1, RD2, US, MUX1_SEL, MUX2_SEL, PC_SEL, RW, WR,
         MEM_ALU_SEL, INST_T_EX, \INST_EX[1] , \INST_EX[0] , \INST_MEM[1] ,
         \INST_MEM[0] ;
  wire   \TMP1E[0] , \TMP2E[0] , \TMP5E[0] , \TMP11M[0] , \TMP12M[0] ,
         \TMP11W[0] , \TMP21W[0] , \TMP12W[0] , \TMP22W[0] , \TMP13W[0] ,
         \TMP23W[0] , \INST_TMP[0] , \INST_TMP1[0] , n177, n178, n179, n181,
         n1, n4, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n180, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202;
  wire   [5:0] OPCODE1;
  wire   [5:0] OPCODE2;
  wire   [5:0] OPCODE3;
  wire   [10:0] FUNC1;
  wire   [1:0] INST;
  wire   [1:0] NEXT_INST;
  wire   [21:0] cw;
  wire   [2:0] TMP3E;
  wire   [3:0] TMP4E;
  wire   [1:0] TMP21M;
  wire   [1:0] TMP22M;
  wire   [1:0] INST1;

  DFFR_X1 \INST_reg[1]  ( .D(NEXT_INST[1]), .CK(CLK), .RN(n20), .Q(INST[1]) );
  DFFR_X1 \INST1_reg[1]  ( .D(INST[1]), .CK(CLK), .RN(n20), .Q(INST1[1]) );
  DFFR_X1 \INST1_reg[0]  ( .D(INST[0]), .CK(CLK), .RN(n20), .Q(INST1[0]) );
  DFFR_X1 \INST2_reg[1]  ( .D(INST1[1]), .CK(CLK), .RN(n20), .Q(INST_EX[1]) );
  DFFR_X1 \INST3_reg[1]  ( .D(INST_EX[1]), .CK(CLK), .RN(n20), .Q(INST_MEM[1])
         );
  NAND3_X1 U198 ( .A1(n178), .A2(n179), .A3(INST[1]), .ZN(n177) );
  DFFR_X1 \INST_reg[0]  ( .D(NEXT_INST[0]), .CK(CLK), .RN(RST), .Q(INST[0]), 
        .QN(n179) );
  DFFR_X1 \INST2_reg[0]  ( .D(INST1[0]), .CK(CLK), .RN(RST), .Q(INST_EX[0]), 
        .QN(n1) );
  OR2_X1 U3 ( .A1(INST[1]), .A2(n179), .ZN(n188) );
  AND2_X1 U4 ( .A1(n29), .A2(n103), .ZN(n10) );
  AND4_X1 U5 ( .A1(n40), .A2(\INST_TMP[0] ), .A3(n39), .A4(n38), .ZN(n15) );
  NAND2_X1 U6 ( .A1(n193), .A2(n199), .ZN(n202) );
  NAND2_X1 U7 ( .A1(n73), .A2(n109), .ZN(n135) );
  OAI221_X1 U8 ( .B1(n27), .B2(n25), .C1(n25), .C2(n133), .A(n185), .ZN(n89)
         );
  NAND2_X1 U9 ( .A1(n157), .A2(n152), .ZN(n199) );
  NOR2_X1 U10 ( .A1(n87), .A2(n22), .ZN(\INST_TMP[0] ) );
  OAI21_X1 U11 ( .B1(n88), .B2(n87), .A(n195), .ZN(cw[19]) );
  NAND4_X1 U12 ( .A1(n130), .A2(n10), .A3(n4), .A4(n33), .ZN(n158) );
  NAND2_X1 U13 ( .A1(n157), .A2(n84), .ZN(n88) );
  NAND2_X1 U14 ( .A1(n35), .A2(n65), .ZN(n123) );
  AND2_X1 U15 ( .A1(n133), .A2(n123), .ZN(n4) );
  NAND2_X1 U16 ( .A1(n146), .A2(n56), .ZN(n196) );
  NAND2_X1 U17 ( .A1(n109), .A2(n67), .ZN(n103) );
  NAND2_X1 U18 ( .A1(n65), .A2(n84), .ZN(n27) );
  NAND2_X1 U19 ( .A1(n153), .A2(n110), .ZN(n185) );
  NAND2_X1 U20 ( .A1(n35), .A2(n144), .ZN(n200) );
  NOR2_X1 U21 ( .A1(n110), .A2(n109), .ZN(n111) );
  AND2_X1 U22 ( .A1(n37), .A2(n151), .ZN(n9) );
  OAI22_X1 U23 ( .A1(n79), .A2(n180), .B1(n85), .B2(n66), .ZN(n159) );
  AOI21_X1 U24 ( .B1(n153), .B2(n26), .A(n89), .ZN(n130) );
  OAI21_X1 U25 ( .B1(n34), .B2(n23), .A(n123), .ZN(n26) );
  OAI21_X1 U26 ( .B1(n182), .B2(n24), .A(n120), .ZN(n110) );
  NAND2_X1 U27 ( .A1(n157), .A2(n15), .ZN(n190) );
  OAI211_X1 U28 ( .C1(n41), .C2(n94), .A(n171), .B(n170), .ZN(n127) );
  NAND2_X1 U29 ( .A1(n35), .A2(n18), .ZN(n133) );
  NAND2_X1 U30 ( .A1(n30), .A2(n122), .ZN(n153) );
  AND4_X1 U31 ( .A1(n50), .A2(n173), .A3(n94), .A4(n49), .ZN(n11) );
  NAND2_X1 U32 ( .A1(n92), .A2(n113), .ZN(n145) );
  NAND2_X1 U33 ( .A1(n138), .A2(n14), .ZN(n172) );
  NAND2_X1 U34 ( .A1(n69), .A2(n80), .ZN(n71) );
  NAND2_X1 U35 ( .A1(n64), .A2(n66), .ZN(n22) );
  NAND2_X1 U36 ( .A1(n68), .A2(n67), .ZN(n80) );
  NAND2_X1 U37 ( .A1(n45), .A2(n44), .ZN(n46) );
  NAND2_X1 U38 ( .A1(n112), .A2(n46), .ZN(n51) );
  NAND2_X1 U39 ( .A1(n21), .A2(n28), .ZN(n81) );
  AND2_X1 U40 ( .A1(n145), .A2(n14), .ZN(n12) );
  OAI22_X1 U41 ( .A1(n172), .A2(n190), .B1(n184), .B2(n188), .ZN(n141) );
  OAI22_X1 U42 ( .A1(n11), .A2(n190), .B1(n130), .B2(n188), .ZN(n131) );
  AND3_X1 U43 ( .A1(n134), .A2(n126), .A3(n125), .ZN(n13) );
  OAI211_X1 U44 ( .C1(n133), .C2(n188), .A(n132), .B(n149), .ZN(cw[6]) );
  OAI211_X1 U45 ( .C1(n151), .C2(n188), .A(n150), .B(n149), .ZN(cw[10]) );
  AND2_X1 U46 ( .A1(n173), .A2(n170), .ZN(n91) );
  NAND2_X1 U47 ( .A1(n152), .A2(n36), .ZN(n151) );
  NOR2_X1 U48 ( .A1(n159), .A2(n71), .ZN(n70) );
  NAND2_X1 U49 ( .A1(n10), .A2(n115), .ZN(n119) );
  AND4_X1 U50 ( .A1(FUNC[2]), .A2(n53), .A3(n43), .A4(n42), .ZN(n14) );
  NAND4_X1 U51 ( .A1(OPCODE[3]), .A2(OPCODE[5]), .A3(OPCODE[1]), .A4(n64), 
        .ZN(n120) );
  AND2_X1 U52 ( .A1(FUNC[5]), .A2(n42), .ZN(n16) );
  AND3_X1 U53 ( .A1(FUNC[5]), .A2(FUNC[4]), .A3(FUNC[3]), .ZN(n17) );
  NAND2_X1 U54 ( .A1(FUNC[1]), .A2(n44), .ZN(n113) );
  NAND2_X1 U55 ( .A1(OPCODE[0]), .A2(n28), .ZN(n180) );
  NAND2_X1 U56 ( .A1(n157), .A2(n78), .ZN(n161) );
  NAND2_X1 U57 ( .A1(OPCODE[0]), .A2(OPCODE[4]), .ZN(n122) );
  NAND2_X1 U58 ( .A1(n45), .A2(FUNC[0]), .ZN(n112) );
  AND2_X1 U59 ( .A1(OPCODE[1]), .A2(OPCODE[3]), .ZN(n18) );
  NAND2_X1 U60 ( .A1(FUNC[1]), .A2(FUNC[0]), .ZN(n92) );
  NAND2_X1 U61 ( .A1(OPCODE[2]), .A2(n66), .ZN(n23) );
  NAND2_X1 U62 ( .A1(OPCODE[1]), .A2(n58), .ZN(n34) );
  NAND2_X1 U63 ( .A1(n57), .A2(OPCODE[3]), .ZN(n24) );
  NAND2_X1 U64 ( .A1(n21), .A2(OPCODE[4]), .ZN(n30) );
  NAND2_X1 U65 ( .A1(OPCODE[2]), .A2(OPCODE[5]), .ZN(n182) );
  NAND2_X1 U66 ( .A1(n177), .A2(n199), .ZN(NEXT_INST[1]) );
  NOR4_X1 U67 ( .A1(OPCODE1[2]), .A2(n181), .A3(OPCODE1[5]), .A4(OPCODE1[3]), 
        .ZN(n178) );
  INV_X1 U68 ( .A(OPCODE1[1]), .ZN(n181) );
  BUF_X2 U69 ( .A(RST), .Z(n20) );
  CLKBUF_X3 U70 ( .A(RST), .Z(n19) );
  INV_X1 U71 ( .A(OPCODE[3]), .ZN(n58) );
  INV_X1 U72 ( .A(OPCODE[0]), .ZN(n21) );
  INV_X1 U73 ( .A(OPCODE[4]), .ZN(n28) );
  INV_X1 U74 ( .A(n81), .ZN(n73) );
  INV_X1 U75 ( .A(OPCODE[1]), .ZN(n57) );
  NAND3_X1 U76 ( .A1(n58), .A2(n73), .A3(n57), .ZN(n87) );
  INV_X1 U77 ( .A(OPCODE[2]), .ZN(n64) );
  INV_X1 U78 ( .A(OPCODE[5]), .ZN(n66) );
  INV_X1 U79 ( .A(n22), .ZN(n35) );
  INV_X1 U80 ( .A(n24), .ZN(n65) );
  INV_X1 U81 ( .A(n23), .ZN(n84) );
  INV_X1 U82 ( .A(n153), .ZN(n25) );
  NAND3_X1 U83 ( .A1(n73), .A2(n84), .A3(n18), .ZN(n29) );
  INV_X1 U84 ( .A(n27), .ZN(n109) );
  INV_X1 U85 ( .A(n180), .ZN(n67) );
  INV_X1 U86 ( .A(n30), .ZN(n31) );
  NAND3_X1 U87 ( .A1(n31), .A2(n84), .A3(n58), .ZN(n184) );
  INV_X1 U88 ( .A(n184), .ZN(n32) );
  INV_X1 U89 ( .A(n135), .ZN(n90) );
  NOR2_X1 U90 ( .A1(n32), .A2(n90), .ZN(n33) );
  INV_X1 U91 ( .A(n158), .ZN(n37) );
  INV_X1 U92 ( .A(n34), .ZN(n144) );
  INV_X1 U93 ( .A(n200), .ZN(n152) );
  NAND2_X1 U94 ( .A1(n122), .A2(n180), .ZN(n36) );
  INV_X1 U95 ( .A(n188), .ZN(n157) );
  INV_X1 U96 ( .A(FUNC[6]), .ZN(n40) );
  INV_X1 U97 ( .A(FUNC[7]), .ZN(n39) );
  NOR3_X1 U98 ( .A1(FUNC[10]), .A2(FUNC[8]), .A3(FUNC[9]), .ZN(n38) );
  INV_X1 U99 ( .A(n190), .ZN(n146) );
  INV_X1 U100 ( .A(FUNC[1]), .ZN(n45) );
  INV_X1 U101 ( .A(n112), .ZN(n164) );
  INV_X1 U102 ( .A(FUNC[0]), .ZN(n44) );
  NOR2_X1 U103 ( .A1(n164), .A2(n145), .ZN(n41) );
  INV_X1 U104 ( .A(FUNC[4]), .ZN(n42) );
  INV_X1 U105 ( .A(FUNC[2]), .ZN(n52) );
  NAND3_X1 U106 ( .A1(FUNC[3]), .A2(n16), .A3(n52), .ZN(n94) );
  INV_X1 U107 ( .A(n113), .ZN(n165) );
  NAND3_X1 U108 ( .A1(n165), .A2(n17), .A3(n52), .ZN(n171) );
  INV_X1 U109 ( .A(n92), .ZN(n163) );
  NAND3_X1 U110 ( .A1(n163), .A2(n17), .A3(n52), .ZN(n170) );
  INV_X1 U111 ( .A(n127), .ZN(n50) );
  NAND3_X1 U112 ( .A1(FUNC[2]), .A2(n17), .A3(n164), .ZN(n173) );
  INV_X1 U113 ( .A(FUNC[3]), .ZN(n53) );
  INV_X1 U114 ( .A(FUNC[5]), .ZN(n43) );
  INV_X1 U115 ( .A(n46), .ZN(n138) );
  NAND3_X1 U116 ( .A1(FUNC[2]), .A2(n138), .A3(n17), .ZN(n167) );
  NAND3_X1 U117 ( .A1(FUNC[2]), .A2(FUNC[3]), .A3(n16), .ZN(n93) );
  INV_X1 U118 ( .A(n93), .ZN(n95) );
  NAND2_X1 U119 ( .A1(n95), .A2(n51), .ZN(n47) );
  NAND2_X1 U120 ( .A1(n167), .A2(n47), .ZN(n48) );
  NOR2_X1 U121 ( .A1(n12), .A2(n48), .ZN(n49) );
  NAND3_X1 U122 ( .A1(FUNC[2]), .A2(n16), .A3(n53), .ZN(n98) );
  INV_X1 U123 ( .A(n98), .ZN(n137) );
  INV_X1 U124 ( .A(n51), .ZN(n97) );
  NAND2_X1 U125 ( .A1(n113), .A2(n97), .ZN(n54) );
  NAND3_X1 U126 ( .A1(n53), .A2(n16), .A3(n52), .ZN(n168) );
  INV_X1 U127 ( .A(n168), .ZN(n129) );
  AOI21_X1 U128 ( .B1(n137), .B2(n54), .A(n129), .ZN(n55) );
  NAND3_X1 U129 ( .A1(n11), .A2(n172), .A3(n55), .ZN(n56) );
  OAI21_X1 U130 ( .B1(n9), .B2(n188), .A(n196), .ZN(cw[0]) );
  NAND2_X1 U131 ( .A1(n15), .A2(n56), .ZN(n155) );
  NAND3_X1 U132 ( .A1(n58), .A2(n67), .A3(n57), .ZN(n85) );
  NAND2_X1 U133 ( .A1(n87), .A2(n85), .ZN(n176) );
  NAND2_X1 U134 ( .A1(OPCODE[5]), .A2(n176), .ZN(n59) );
  NAND2_X1 U135 ( .A1(n155), .A2(n59), .ZN(n62) );
  NOR2_X1 U136 ( .A1(n66), .A2(OPCODE[2]), .ZN(n60) );
  NAND3_X1 U137 ( .A1(n144), .A2(n67), .A3(n60), .ZN(n69) );
  NAND2_X1 U138 ( .A1(n9), .A2(n69), .ZN(n61) );
  OAI21_X1 U139 ( .B1(n62), .B2(n61), .A(n157), .ZN(n63) );
  INV_X1 U140 ( .A(n63), .ZN(cw[1]) );
  NAND3_X1 U141 ( .A1(OPCODE[5]), .A2(n65), .A3(n64), .ZN(n79) );
  INV_X1 U142 ( .A(n120), .ZN(n68) );
  NOR2_X1 U143 ( .A1(n70), .A2(n188), .ZN(cw[3]) );
  INV_X1 U144 ( .A(n71), .ZN(n77) );
  INV_X1 U145 ( .A(n79), .ZN(n72) );
  NAND2_X1 U146 ( .A1(n73), .A2(n72), .ZN(n76) );
  INV_X1 U147 ( .A(n87), .ZN(n74) );
  NAND2_X1 U148 ( .A1(OPCODE[5]), .A2(n74), .ZN(n75) );
  NAND3_X1 U149 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n78) );
  INV_X1 U150 ( .A(n161), .ZN(cw[2]) );
  NAND2_X1 U151 ( .A1(n80), .A2(n79), .ZN(n83) );
  NAND2_X1 U152 ( .A1(n81), .A2(n180), .ZN(n82) );
  NAND3_X1 U153 ( .A1(n157), .A2(n83), .A3(n82), .ZN(n192) );
  INV_X1 U154 ( .A(n192), .ZN(cw[4]) );
  INV_X1 U155 ( .A(n85), .ZN(n86) );
  INV_X1 U156 ( .A(n88), .ZN(n143) );
  NAND2_X1 U157 ( .A1(n86), .A2(n143), .ZN(n195) );
  INV_X1 U158 ( .A(cw[19]), .ZN(n193) );
  NOR2_X1 U159 ( .A1(n90), .A2(n89), .ZN(n107) );
  OAI221_X1 U160 ( .B1(n93), .B2(n112), .C1(n92), .C2(n94), .A(n91), .ZN(n108)
         );
  INV_X1 U161 ( .A(n108), .ZN(n102) );
  NOR2_X1 U162 ( .A1(n113), .A2(n94), .ZN(n100) );
  NAND2_X1 U163 ( .A1(n138), .A2(n95), .ZN(n96) );
  OAI21_X1 U164 ( .B1(n98), .B2(n97), .A(n96), .ZN(n99) );
  NOR2_X1 U165 ( .A1(n100), .A2(n99), .ZN(n101) );
  NAND4_X1 U166 ( .A1(n171), .A2(n102), .A3(n167), .A4(n101), .ZN(n105) );
  INV_X1 U167 ( .A(n103), .ZN(n104) );
  AOI21_X1 U168 ( .B1(n15), .B2(n105), .A(n104), .ZN(n106) );
  AOI21_X1 U169 ( .B1(n107), .B2(n106), .A(n188), .ZN(cw[9]) );
  NAND2_X1 U170 ( .A1(n146), .A2(n108), .ZN(n118) );
  AOI21_X1 U171 ( .B1(n133), .B2(n111), .A(n122), .ZN(n116) );
  NAND2_X1 U172 ( .A1(n113), .A2(n112), .ZN(n114) );
  NAND3_X1 U173 ( .A1(n15), .A2(n137), .A3(n114), .ZN(n115) );
  OAI21_X1 U174 ( .B1(n116), .B2(n119), .A(n157), .ZN(n117) );
  NAND2_X1 U175 ( .A1(n118), .A2(n117), .ZN(cw[8]) );
  INV_X1 U176 ( .A(n119), .ZN(n134) );
  NAND2_X1 U177 ( .A1(n133), .A2(n120), .ZN(n121) );
  NAND2_X1 U178 ( .A1(n153), .A2(n121), .ZN(n126) );
  INV_X1 U179 ( .A(n122), .ZN(n142) );
  INV_X1 U180 ( .A(n123), .ZN(n124) );
  NAND2_X1 U181 ( .A1(n142), .A2(n124), .ZN(n125) );
  NAND2_X1 U182 ( .A1(n146), .A2(n127), .ZN(n128) );
  OAI21_X1 U183 ( .B1(n13), .B2(n188), .A(n128), .ZN(cw[7]) );
  NAND3_X1 U184 ( .A1(n129), .A2(n145), .A3(n146), .ZN(n132) );
  INV_X1 U185 ( .A(n131), .ZN(n149) );
  NAND3_X1 U186 ( .A1(n135), .A2(n134), .A3(n151), .ZN(n136) );
  NAND2_X1 U187 ( .A1(n157), .A2(n136), .ZN(n140) );
  NAND3_X1 U188 ( .A1(n146), .A2(n138), .A3(n137), .ZN(n139) );
  NAND2_X1 U189 ( .A1(n140), .A2(n139), .ZN(cw[12]) );
  INV_X1 U190 ( .A(n141), .ZN(n150) );
  NAND3_X1 U191 ( .A1(n144), .A2(n143), .A3(n142), .ZN(n148) );
  NAND3_X1 U192 ( .A1(n146), .A2(n14), .A3(n145), .ZN(n147) );
  NAND3_X1 U193 ( .A1(n150), .A2(n148), .A3(n147), .ZN(cw[11]) );
  NAND2_X1 U194 ( .A1(n153), .A2(n152), .ZN(n154) );
  NAND2_X1 U195 ( .A1(n155), .A2(n154), .ZN(n156) );
  NAND2_X1 U196 ( .A1(n157), .A2(n156), .ZN(n162) );
  INV_X1 U197 ( .A(n162), .ZN(cw[13]) );
  OAI21_X1 U199 ( .B1(n159), .B2(n158), .A(n157), .ZN(n160) );
  NAND2_X1 U200 ( .A1(n161), .A2(n160), .ZN(cw[20]) );
  INV_X1 U201 ( .A(cw[20]), .ZN(n198) );
  NAND2_X1 U202 ( .A1(n198), .A2(n162), .ZN(cw[14]) );
  NOR2_X1 U203 ( .A1(n164), .A2(n163), .ZN(n169) );
  NAND2_X1 U204 ( .A1(n165), .A2(n14), .ZN(n166) );
  OAI211_X1 U205 ( .C1(n169), .C2(n168), .A(n167), .B(n166), .ZN(n175) );
  NAND4_X1 U206 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .ZN(n174) );
  NOR2_X1 U207 ( .A1(n175), .A2(n174), .ZN(n191) );
  INV_X1 U208 ( .A(n176), .ZN(n183) );
  OAI22_X1 U209 ( .A1(n183), .A2(n182), .B1(n4), .B2(n180), .ZN(n187) );
  NAND2_X1 U210 ( .A1(n185), .A2(n184), .ZN(n186) );
  NOR2_X1 U211 ( .A1(n187), .A2(n186), .ZN(n189) );
  OAI22_X1 U212 ( .A1(n191), .A2(n190), .B1(n189), .B2(n188), .ZN(cw[15]) );
  NAND2_X1 U213 ( .A1(n196), .A2(n192), .ZN(cw[16]) );
  INV_X1 U214 ( .A(cw[14]), .ZN(n194) );
  NAND2_X1 U215 ( .A1(n194), .A2(n193), .ZN(cw[17]) );
  INV_X1 U216 ( .A(n195), .ZN(cw[18]) );
  INV_X1 U217 ( .A(n199), .ZN(cw[21]) );
  INV_X1 U218 ( .A(n202), .ZN(n197) );
  NAND3_X1 U219 ( .A1(n198), .A2(n197), .A3(n196), .ZN(STALL) );
  NOR2_X1 U220 ( .A1(n200), .A2(n179), .ZN(n201) );
  OAI22_X1 U221 ( .A1(n178), .A2(INST[0]), .B1(n201), .B2(INST[1]), .ZN(
        NEXT_INST[0]) );
  FD_NB6_3 OPPP1 ( .CK(CLK), .RESET(n19), .D(OPCODE), .Q(OPCODE1) );
  FD_NB6_2 OPPP2 ( .CK(CLK), .RESET(n19), .D(OPCODE1), .Q(OPCODE2) );
  FD_NB6_1 OPPP3 ( .CK(CLK), .RESET(n19), .D(OPCODE2), .Q(OPCODE3) );
  FD_NB6_0 OPPP4 ( .CK(CLK), .RESET(n19), .D(OPCODE3) );
  FD_NB11_1 FUNPP1 ( .CK(CLK), .RESET(n19), .D(FUNC), .Q(FUNC1) );
  FD_NB11_0 FUNPP2 ( .CK(CLK), .RESET(n19), .D(FUNC1) );
  FD_NB1_22 pipe1_JMP ( .CK(CLK), .RESET(n20), .D(cw[21]), .Q(JMP) );
  FD_NB1_21 pipe1_RI ( .CK(CLK), .RESET(n20), .D(cw[20]), .Q(RI) );
  FD_NB2_3 pipe1_BR ( .CK(CLK), .RESET(n20), .D(cw[19:18]), .Q(BR_TYPE) );
  FD_NB1_20 pipe1_RD1 ( .CK(CLK), .RESET(n20), .D(cw[17]), .Q(RD1) );
  FD_NB1_19 pipe1_RD2 ( .CK(CLK), .RESET(n20), .D(cw[16]), .Q(RD2) );
  FD_NB1_18 pipe1_US ( .CK(CLK), .RESET(n20), .D(cw[15]), .Q(US) );
  FD_NB1_17 pipe1_MX1 ( .CK(CLK), .RESET(n20), .D(cw[14]), .Q(\TMP1E[0] ) );
  FD_NB1_16 pipe1_MX2 ( .CK(CLK), .RESET(n20), .D(cw[13]), .Q(\TMP2E[0] ) );
  FD_NB3_1 pipe1_UN ( .CK(CLK), .RESET(n20), .D(cw[12:10]), .Q(TMP3E) );
  FD_NB4_1 pipe1_OP ( .CK(CLK), .RESET(n19), .D(cw[9:6]), .Q(TMP4E) );
  FD_NB1_15 pipe1_PC ( .CK(CLK), .RESET(n20), .D(n202), .Q(\TMP5E[0] ) );
  FD_NB1_14 pipe2_MX1 ( .CK(CLK), .RESET(n20), .D(\TMP1E[0] ), .Q(MUX1_SEL) );
  FD_NB1_13 pipe2_MX2 ( .CK(CLK), .RESET(n20), .D(\TMP2E[0] ), .Q(MUX2_SEL) );
  FD_NB3_0 pipe2_UN ( .CK(CLK), .RESET(n20), .D(TMP3E), .Q(UN_SEL) );
  FD_NB4_0 pipe2_OP ( .CK(CLK), .RESET(n19), .D(TMP4E), .Q(OP_SEL) );
  FD_NB1_12 pipe2_PC ( .CK(CLK), .RESET(n20), .D(\TMP5E[0] ), .Q(PC_SEL) );
  FD_NB1_11 pipe1_RW ( .CK(CLK), .RESET(n20), .D(cw[4]), .Q(\TMP11M[0] ) );
  FD_NB2_2 pipe1_DT ( .CK(CLK), .RESET(n20), .D(cw[3:2]), .Q(TMP21M) );
  FD_NB1_10 pipe2_RW ( .CK(CLK), .RESET(n20), .D(\TMP11M[0] ), .Q(\TMP12M[0] )
         );
  FD_NB2_1 pipe2_DT ( .CK(CLK), .RESET(n20), .D(TMP21M), .Q(TMP22M) );
  FD_NB1_9 pipe3_RW ( .CK(CLK), .RESET(n20), .D(\TMP12M[0] ), .Q(RW) );
  FD_NB2_0 pipe3_DT ( .CK(CLK), .RESET(n20), .D(TMP22M), .Q(D_TYPE) );
  FD_INJ_NB1_2 pipe1_WR ( .CK(CLK), .RESET(n20), .INJ_ZERO(FLUSH), .D(cw[1]), 
        .Q(\TMP11W[0] ) );
  FD_NB1_8 pipe1_MM ( .CK(CLK), .RESET(n20), .D(cw[0]), .Q(\TMP21W[0] ) );
  FD_INJ_NB1_1 pipe2_WR ( .CK(CLK), .RESET(FLUSH), .INJ_ZERO(n20), .D(
        \TMP11W[0] ), .Q(\TMP12W[0] ) );
  FD_NB1_7 pipe2_MM ( .CK(CLK), .RESET(n20), .D(\TMP21W[0] ), .Q(\TMP22W[0] )
         );
  FD_NB1_6 pipe3_WR ( .CK(CLK), .RESET(n20), .D(\TMP12W[0] ), .Q(\TMP13W[0] )
         );
  FD_NB1_5 pipe3_MM ( .CK(CLK), .RESET(n20), .D(\TMP22W[0] ), .Q(\TMP23W[0] )
         );
  FD_NB1_4 pipe4_WR ( .CK(CLK), .RESET(n20), .D(\TMP13W[0] ), .Q(WR) );
  FD_NB1_3 pipe4_MM ( .CK(CLK), .RESET(n20), .D(\TMP23W[0] ), .Q(MEM_ALU_SEL)
         );
  FD_NB1_2 pipe1_INST ( .CK(CLK), .RESET(n20), .D(\INST_TMP[0] ), .Q(
        \INST_TMP1[0] ) );
  FD_NB1_1 pipe2_INST ( .CK(CLK), .RESET(n20), .D(\INST_TMP1[0] ), .Q(
        INST_T_EX) );
  SDFFR_X1 \INST3_reg[0]  ( .D(1'b1), .SI(1'b0), .SE(n1), .CK(CLK), .RN(n20), 
        .Q(INST_MEM[0]) );
endmodule


module DATAPATH_NB32_LS5_OPC6_FN11_0 ( CLK, STALL, RST, .INST_EX({\INST_EX[1] , 
        \INST_EX[0] }), .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }), INST_T_EX, 
        JMP, RI, RD1, RD2, WR, PC_SEL, MEM_ALU_SEL, US, MUX1_SEL, MUX2_SEL, 
        BR_TYPE, UN_SEL, OP_SEL, IRAM_OUT, EXT_MEM_IN, FLUSH, US_MEM, HAZARD, 
        EXT_MEM_ADD, EXT_MEM_DATA, CURR_PC, FUNC, OP_CODE );
  input [1:0] BR_TYPE;
  input [2:0] UN_SEL;
  input [3:0] OP_SEL;
  input [31:0] IRAM_OUT;
  input [31:0] EXT_MEM_IN;
  output [4:0] EXT_MEM_ADD;
  output [31:0] EXT_MEM_DATA;
  output [31:0] CURR_PC;
  output [10:0] FUNC;
  output [5:0] OP_CODE;
  input CLK, STALL, RST, \INST_EX[1] , \INST_EX[0] , \INST_MEM[1] ,
         \INST_MEM[0] , INST_T_EX, JMP, RI, RD1, RD2, WR, PC_SEL, MEM_ALU_SEL,
         US, MUX1_SEL, MUX2_SEL;
  output FLUSH, US_MEM, HAZARD;
  wire   n13, US_TO_EX, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12;
  wire   [1:0] MISS_HIT;
  wire   [31:0] TEMP_PC;
  wire   [31:0] NPC;
  wire   [25:0] INST;
  wire   [31:0] DATA_WB;
  wire   [4:0] DEST_FROM_WRBU;
  wire   [31:0] A;
  wire   [31:0] B;
  wire   [31:0] C;
  wire   [31:0] D;
  wire   [4:0] RT;
  wire   [4:0] RS;
  wire   [4:0] DEST_FROM_DECU;
  wire   [1:0] FW_MUX1_SEL;
  wire   [1:0] FW_MUX2_SEL;
  wire   [31:5] ALU_OUT;
  wire   [4:0] DEST_FROM_EXEU;
  wire   [31:0] ALU_TO_WB;
  wire   [31:0] TMP_MEM;
  wire   [4:0] DEST_FROM_MEMU;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5;

  CLKBUF_X3 U1 ( .A(n13), .Z(FLUSH) );
  CLKBUF_X1 U2 ( .A(DEST_FROM_MEMU[4]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(DEST_FROM_MEMU[1]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(DEST_FROM_MEMU[2]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(DEST_FROM_EXEU[0]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(DEST_FROM_MEMU[3]), .Z(n5) );
  INV_X1 U7 ( .A(RST), .ZN(n12) );
  CLKBUF_X1 U8 ( .A(DEST_FROM_EXEU[2]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(DEST_FROM_EXEU[3]), .Z(n7) );
  CLKBUF_X1 U10 ( .A(DEST_FROM_EXEU[4]), .Z(n8) );
  CLKBUF_X1 U11 ( .A(DEST_FROM_EXEU[1]), .Z(n9) );
  CLKBUF_X1 U12 ( .A(DEST_FROM_MEMU[0]), .Z(n10) );
  AOI21_X1 U13 ( .B1(MISS_HIT[1]), .B2(MISS_HIT[0]), .A(n12), .ZN(n13) );
  FETCH_UNIT_NB32_LS5_0 ife_unit ( .CLK(CLK), .STALL(STALL), .RST(RST), 
        .RST_DEC(RST), .PC_SEL(PC_SEL), .JB_INST(TEMP_PC), .IRAM_OUT(IRAM_OUT), 
        .FUNC(FUNC), .OPCODE(OP_CODE), .CURR_PC(CURR_PC), .NPC(NPC), 
        .INST_OUT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, INST}), .MISS_HIT(
        MISS_HIT) );
  DECODE_UNIT_NB32_LS5_0 dec_unit ( .CLK(CLK), .RST(RST), .FLUSH(FLUSH), 
        .DATAIN(DATA_WB), .IMM1(INST), .IMM2(NPC), .BR_TYPE(BR_TYPE), .JMP(JMP), .RI(RI), .US(US), .RD1(RD1), .RD2(RD2), .WR(WR), .ADD_WR(DEST_FROM_WRBU), 
        .ADD_RD1(INST[25:21]), .ADD_RD2(INST[20:16]), .DEST_IN(INST[15:11]), 
        .HAZARD(HAZARD), .US_TO_EX(US_TO_EX), .A(A), .B(B), .C(C), .D(D), .RT(
        RT), .RS(RS), .DEST_OUT(DEST_FROM_DECU) );
  EXECUTION_UNIT_NB32_LS5_0 exe_unit ( .FW_MUX1_SEL(FW_MUX1_SEL), 
        .FW_MUX2_SEL(FW_MUX2_SEL), .FW_EX({ALU_OUT, EXT_MEM_ADD}), .FW_MEM(
        DATA_WB), .A(A), .B(B), .C(C), .D(D), .DEST_IN(DEST_FROM_DECU), .CLK(
        CLK), .RST(RST), .US(US_TO_EX), .MUX1_SEL(MUX1_SEL), .MUX2_SEL(
        MUX2_SEL), .UN_SEL(UN_SEL), .OP_SEL(OP_SEL), .US_MEM(US_MEM), 
        .TEMP_PC(TEMP_PC), .ALU_OUT({ALU_OUT, EXT_MEM_ADD}), .IMM_OUT(
        EXT_MEM_DATA), .DEST_OUT(DEST_FROM_EXEU) );
  MEMORY_UNIT_NB32_LS5_0 mem_unit ( .CLK(CLK), .RST(RST), .DEST_IN({n8, n7, n6, 
        n9, n4}), .FROM_MEM(EXT_MEM_IN), .FROM_ALU({ALU_OUT, EXT_MEM_ADD}), 
        .ALU_OUT(ALU_TO_WB), .MEM_OUT(TMP_MEM), .DEST_OUT(DEST_FROM_MEMU) );
  WRITE_BACK_UNIT_NB32_LS5_0 wrb_unit ( .MEM_ALU_SEL(MEM_ALU_SEL), .DEST_IN({
        n1, n5, n3, n2, n10}), .FROM_ALU(ALU_TO_WB), .FROM_MEM(TMP_MEM), 
        .DATA_OUT(DATA_WB), .DEST_OUT(DEST_FROM_WRBU) );
  FOREWARD_UNIT_NB32_LS5_0 fw_unit ( .INST_EX({\INST_EX[1] , \INST_EX[0] }), 
        .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }), .INST_T_EX(INST_T_EX), 
        .Rs_EX(RS), .Rt_EX(RT), .Rd_MEM(DEST_FROM_EXEU), .Rd_WB(DEST_FROM_MEMU), .CTL_MUX1(FW_MUX1_SEL), .CTL_MUX2(FW_MUX2_SEL) );
endmodule


module DLX ( CLK, RST, D_TYPE, EXT_MEM_IN, IRAM_OUT, RW, US_MEM, IRAM_ADD, 
        EXT_MEM_ADD, EXT_MEM_DATA );
  output [1:0] D_TYPE;
  input [31:0] EXT_MEM_IN;
  input [31:0] IRAM_OUT;
  output [31:0] IRAM_ADD;
  output [4:0] EXT_MEM_ADD;
  output [31:0] EXT_MEM_DATA;
  input CLK, RST;
  output RW, US_MEM;
  wire   STALL, INST_T_EX, JMP, RI, RD1, RD2, WR, PC_SEL, MEM_ALU_SEL, US,
         MUX1_SEL, MUX2_SEL, FLUSH;
  wire   [1:0] INST_EX;
  wire   [1:0] INST_MEM;
  wire   [1:0] BR_TYPE;
  wire   [2:0] UN_SEL;
  wire   [3:0] OP_SEL;
  wire   [10:0] FUNC;
  wire   [5:0] OPCODE;

  DATAPATH_NB32_LS5_OPC6_FN11_0 dp ( .CLK(CLK), .STALL(STALL), .RST(RST), 
        .INST_EX(INST_EX), .INST_MEM(INST_MEM), .INST_T_EX(INST_T_EX), .JMP(
        JMP), .RI(RI), .RD1(RD1), .RD2(RD2), .WR(WR), .PC_SEL(PC_SEL), 
        .MEM_ALU_SEL(MEM_ALU_SEL), .US(US), .MUX1_SEL(MUX1_SEL), .MUX2_SEL(
        MUX2_SEL), .BR_TYPE(BR_TYPE), .UN_SEL(UN_SEL), .OP_SEL(OP_SEL), 
        .IRAM_OUT(IRAM_OUT), .EXT_MEM_IN(EXT_MEM_IN), .FLUSH(FLUSH), .US_MEM(
        US_MEM), .EXT_MEM_ADD(EXT_MEM_ADD), .EXT_MEM_DATA(EXT_MEM_DATA), 
        .CURR_PC(IRAM_ADD), .FUNC(FUNC), .OP_CODE(OPCODE) );
  DLX_CU_0 cu ( .CLK(CLK), .RST(RST), .OPCODE(OPCODE), .FUNC(FUNC), .FLUSH(
        FLUSH), .STALL(STALL), .JMP(JMP), .RI(RI), .BR_TYPE(BR_TYPE), .RD1(RD1), .RD2(RD2), .US(US), .MUX1_SEL(MUX1_SEL), .MUX2_SEL(MUX2_SEL), .UN_SEL(UN_SEL), .OP_SEL(OP_SEL), .PC_SEL(PC_SEL), .RW(RW), .D_TYPE(D_TYPE), .WR(WR), 
        .MEM_ALU_SEL(MEM_ALU_SEL), .INST_T_EX(INST_T_EX), .INST_EX(INST_EX), 
        .INST_MEM(INST_MEM) );
endmodule

