
module carry_sel_bk_NB4_49 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  NOR2_X1 U7 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  OAI22_X1 U9 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U10 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U11 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U12 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U16 ( .A(B[1]), .ZN(n56) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_32 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n46), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(B[1]), .ZN(n56) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n46), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n46), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n46), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U14 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U17 ( .A(Ci), .ZN(n46) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_33 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  INV_X1 U16 ( .A(B[1]), .ZN(n56) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_25 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  INV_X1 U3 ( .A(B[1]), .ZN(n56) );
  NAND2_X1 U4 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U5 ( .A(n53), .ZN(n48) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  NOR2_X1 U11 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  OAI22_X1 U12 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_17 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U3 ( .A(n53), .ZN(n48) );
  OAI22_X1 U4 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  INV_X1 U6 ( .A(Ci), .ZN(n68) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  INV_X1 U16 ( .A(B[1]), .ZN(n56) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_34 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  INV_X1 U16 ( .A(B[1]), .ZN(n56) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_26 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  INV_X1 U3 ( .A(B[1]), .ZN(n56) );
  NAND2_X1 U4 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U5 ( .A(n53), .ZN(n48) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  NOR2_X1 U11 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  OAI22_X1 U12 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_23 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  NOR2_X1 U10 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NAND2_X1 U13 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U16 ( .A(B[1]), .ZN(n56) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_15 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  INV_X1 U16 ( .A(B[1]), .ZN(n56) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_58 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NOR2_X1 U14 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U17 ( .A(B[1]), .ZN(n56) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_57 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  AOI22_X1 U12 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U17 ( .A(B[1]), .ZN(n56) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_14 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U4 ( .A(n53), .ZN(n48) );
  OAI22_X1 U5 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NOR2_X1 U9 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U10 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  INV_X1 U11 ( .A(B[1]), .ZN(n56) );
  OAI22_X1 U12 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U13 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U14 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U15 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_61 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  INV_X1 U3 ( .A(A[1]), .ZN(n56) );
  NAND2_X1 U4 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U5 ( .A(n52), .ZN(n47) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(B[1]), .ZN(n55) );
endmodule


module carry_sel_bk_NB4_54 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U3 ( .A(n52), .ZN(n47) );
  INV_X1 U4 ( .A(Ci), .ZN(n68) );
  NOR2_X1 U5 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U9 ( .A(A[1]), .ZN(n56) );
  OAI22_X1 U10 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U12 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U13 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U14 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U15 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(B[1]), .ZN(n55) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_53 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  NOR2_X1 U5 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U9 ( .A(A[1]), .ZN(n56) );
  OAI22_X1 U10 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U12 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U13 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U14 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U15 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(B[1]), .ZN(n55) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_46 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U16 ( .A(A[1]), .ZN(n56) );
  INV_X1 U17 ( .A(B[1]), .ZN(n55) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_45 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U16 ( .A(A[1]), .ZN(n56) );
  INV_X1 U17 ( .A(B[1]), .ZN(n55) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_44 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  OAI22_X1 U7 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U9 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U16 ( .A(A[1]), .ZN(n56) );
  INV_X1 U17 ( .A(B[1]), .ZN(n55) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_38 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_37 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_36 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_29 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_28 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_21 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_20 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_55 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U3 ( .A(n52), .ZN(n47) );
  INV_X1 U4 ( .A(Ci), .ZN(n68) );
  NOR2_X1 U5 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U9 ( .A(A[1]), .ZN(n56) );
  OAI22_X1 U10 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U12 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U13 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U14 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U15 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(B[1]), .ZN(n55) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_31 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  INV_X1 U3 ( .A(B[1]), .ZN(n56) );
  NAND2_X1 U4 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U5 ( .A(n53), .ZN(n48) );
  OAI22_X1 U6 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_27 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_19 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  NAND2_X1 U3 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U4 ( .A(n52), .ZN(n47) );
  OAI22_X1 U5 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U7 ( .A(B[1]), .ZN(n55) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  INV_X1 U3 ( .A(B[1]), .ZN(n55) );
  NAND2_X1 U4 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U5 ( .A(n52), .ZN(n47) );
  OAI22_X1 U6 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U7 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  OAI22_X1 U8 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  OAI22_X1 U10 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NOR2_X1 U14 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  NOR2_X1 U15 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U17 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
endmodule


module carry_sel_bk_NB4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n54), .B(n50), .Z(n51) );
  XOR2_X1 U25 ( .A(n53), .B(n50), .Z(n52) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n50) );
  XOR2_X1 U27 ( .A(n68), .B(n49), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  OAI22_X1 U3 ( .A1(n47), .A2(n56), .B1(n55), .B2(n54), .ZN(n63) );
  OAI22_X1 U4 ( .A1(n47), .A2(n56), .B1(n53), .B2(n55), .ZN(n60) );
  INV_X1 U5 ( .A(B[1]), .ZN(n56) );
  NAND2_X1 U6 ( .A1(n48), .A2(n54), .ZN(n49) );
  INV_X1 U7 ( .A(n53), .ZN(n48) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n53) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  AOI22_X1 U10 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U13 ( .A1(B[0]), .A2(A[0]), .ZN(n54) );
  OR2_X1 U14 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  OAI22_X1 U15 ( .A1(n68), .A2(n52), .B1(Ci), .B2(n51), .ZN(S[1]) );
  OAI22_X1 U16 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  OAI22_X1 U17 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  OAI22_X1 U3 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U4 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U5 ( .A(B[1]), .ZN(n55) );
  NAND2_X1 U6 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U7 ( .A(n52), .ZN(n47) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  AOI22_X1 U10 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U13 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U14 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U15 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  OAI22_X1 U16 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
  OAI22_X1 U17 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U18 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
endmodule


module carry_sel_bk_NB4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  XOR2_X1 U19 ( .A(n65), .B(n64), .Z(n66) );
  XOR2_X1 U20 ( .A(n61), .B(n64), .Z(n67) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n64) );
  XOR2_X1 U22 ( .A(n63), .B(n57), .Z(n58) );
  XOR2_X1 U23 ( .A(n60), .B(n57), .Z(n59) );
  XOR2_X1 U24 ( .A(n53), .B(n49), .Z(n50) );
  XOR2_X1 U25 ( .A(n52), .B(n49), .Z(n51) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n49) );
  XOR2_X1 U27 ( .A(n68), .B(n48), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n68) );
  OAI22_X1 U3 ( .A1(n56), .A2(n55), .B1(n54), .B2(n53), .ZN(n63) );
  OAI22_X1 U4 ( .A1(n56), .A2(n55), .B1(n52), .B2(n54), .ZN(n60) );
  INV_X1 U5 ( .A(B[1]), .ZN(n55) );
  NAND2_X1 U6 ( .A1(n47), .A2(n53), .ZN(n48) );
  INV_X1 U7 ( .A(n52), .ZN(n47) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(B[2]), .B1(n60), .B2(n62), .ZN(n61) );
  NOR2_X1 U9 ( .A1(A[0]), .A2(B[0]), .ZN(n52) );
  AOI22_X1 U10 ( .A1(n63), .A2(n62), .B1(B[2]), .B2(A[2]), .ZN(n65) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n57) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U13 ( .A1(B[0]), .A2(A[0]), .ZN(n53) );
  INV_X1 U14 ( .A(A[1]), .ZN(n56) );
  OR2_X1 U15 ( .A1(B[2]), .A2(A[2]), .ZN(n62) );
  OAI22_X1 U16 ( .A1(n68), .A2(n51), .B1(Ci), .B2(n50), .ZN(S[1]) );
  OAI22_X1 U17 ( .A1(n68), .A2(n59), .B1(Ci), .B2(n58), .ZN(S[2]) );
  OAI22_X1 U18 ( .A1(n68), .A2(n67), .B1(Ci), .B2(n66), .ZN(S[3]) );
endmodule


module G_78 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n4;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gij) );
endmodule


module G_80 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n4;

  AOI21_X1 U1 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Gij) );
endmodule


module G_75 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n4) );
endmodule


module G_74 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n4) );
endmodule


module G_73 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n4) );
endmodule


module G_72 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_71 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_70 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_69 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_68 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_67 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_66 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_65 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_64 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_63 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_62 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_61 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_60 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_59 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_58 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_57 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_56 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_55 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_54 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_53 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_52 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_51 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_50 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_49 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_48 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_47 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_46 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_45 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_44 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_43 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_42 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_41 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_40 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_39 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_38 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_37 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_36 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_35 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_34 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_33 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_32 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_31 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_30 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_29 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_28 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_27 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_26 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_25 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_24 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_23 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_22 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_21 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_20 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_19 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_18 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_17 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_16 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_15 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_14 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_13 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_12 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_11 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_10 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_9 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_8 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_7 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_6 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_5 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_4 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_3 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_2 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module G_1 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module blockPG_231 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n4) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_242 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
endmodule


module blockPG_240 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
endmodule


module blockPG_239 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gij) );
endmodule


module blockPG_238 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  INV_X1 U2 ( .A(n5), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_236 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_235 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_234 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
endmodule


module blockPG_233 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
endmodule


module blockPG_232 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_228 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gij) );
endmodule


module blockPG_226 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
endmodule


module blockPG_224 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_223 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_221 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gij) );
endmodule


module blockPG_227 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  INV_X1 U3 ( .A(n5), .ZN(Gij) );
endmodule


module blockPG_225 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_220 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_217 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n5;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n5), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n5) );
endmodule


module blockPG_48 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_229 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_222 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_216 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_215 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_214 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_213 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_212 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_210 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_209 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_208 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_205 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_204 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_200 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_199 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_198 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_197 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_196 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_195 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_193 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_189 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_188 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_187 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_186 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_185 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_183 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_182 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_181 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_178 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_177 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_173 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_172 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_171 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_170 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_169 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_168 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_166 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_162 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_161 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_160 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_159 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_158 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_156 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_155 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_154 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_151 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_150 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_146 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_145 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_144 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_143 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_142 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_141 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_139 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_135 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_134 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_133 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_132 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_131 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_129 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_128 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_127 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_124 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_123 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_119 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_118 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_117 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_116 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_115 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_114 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_112 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_108 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_107 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_106 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_105 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_102 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_101 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_100 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_97 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_96 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_92 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_91 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_90 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_89 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_88 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_87 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_85 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_81 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_80 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_79 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_78 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_77 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_75 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_74 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_73 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_70 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n3), .ZN(Gij) );
endmodule


module blockPG_69 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_65 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_64 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_63 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_62 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_61 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_60 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_58 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_54 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_53 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_52 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_51 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_50 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_47 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_46 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_43 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_42 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_38 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_37 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_36 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_35 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_34 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_33 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_31 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_27 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_26 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_25 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_24 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_23 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_20 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_19 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_16 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_15 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_11 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_10 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_9 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_8 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_7 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_6 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_4 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_218 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_211 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_207 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_206 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_203 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_202 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_192 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_184 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_180 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_179 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_176 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_175 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_165 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_157 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_153 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_152 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_149 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_148 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_138 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_130 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_126 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_125 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_122 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_121 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_111 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_103 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_99 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_98 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_95 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_94 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_84 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_76 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_72 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_71 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_68 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_67 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_57 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_49 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_45 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_44 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_41 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_40 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_30 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_21 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_18 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_17 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_14 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_13 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_3 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_194 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_191 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_190 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_174 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_167 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_164 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_163 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_147 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_140 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_137 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_136 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_120 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_113 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_110 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_109 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_93 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_86 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_83 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_82 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_66 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_59 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_56 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_55 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_39 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_32 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_29 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_28 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_22 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_12 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_5 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_2 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module blockPG_1 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module pg_net_286 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_284 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_283 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_282 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_279 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_278 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_275 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_274 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_273 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_271 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_270 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_267 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_266 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_262 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_281 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_280 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_277 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_276 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_272 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_269 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_268 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_265 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_264 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_261 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_259 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_258 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_257 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_256 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_255 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_254 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_253 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_252 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_251 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_250 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_249 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_248 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_247 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_246 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_245 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_244 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_243 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_242 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_241 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_240 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_239 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_238 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_237 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_236 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_235 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_234 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_233 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_232 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_231 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_230 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_229 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_228 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_227 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_226 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_225 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_224 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_223 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_222 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_221 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_220 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_219 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_218 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_217 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_216 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_215 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_214 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_213 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_212 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_211 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_210 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_209 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_208 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_207 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_206 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_205 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_204 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_203 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_202 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_201 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_200 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_199 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_198 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_197 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_196 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_195 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_194 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_193 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_192 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_191 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_190 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_189 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_188 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_187 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_186 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_185 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_184 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_183 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_182 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_181 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_180 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_179 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_178 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_177 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_176 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_175 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_174 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_173 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_172 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_171 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_170 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_169 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_168 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_167 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_166 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_165 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_164 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_163 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_162 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_161 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_160 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_159 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_158 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_157 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_156 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_155 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_154 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_153 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_152 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_151 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_150 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_149 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_148 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_147 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_146 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_145 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_144 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_143 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_142 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_141 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_140 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_139 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_138 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_137 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_136 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_135 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_134 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_133 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_132 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_131 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_130 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_129 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_128 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_127 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_126 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_125 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_124 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_123 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_122 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_121 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_120 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_119 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_118 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_117 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_116 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_115 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_114 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_113 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_112 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_111 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_110 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_109 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_108 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_107 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_106 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_105 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_104 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_103 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_102 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_101 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_100 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_99 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_98 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_97 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_96 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_95 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_94 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_93 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_92 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_91 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_90 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_89 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_88 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_87 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_86 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_85 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_84 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_83 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_82 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_81 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_80 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_79 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_78 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_77 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_76 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_75 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_74 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_73 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_72 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_71 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_70 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_69 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_68 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_67 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_66 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_65 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_64 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_63 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_62 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_61 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_60 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_59 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_58 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_57 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_56 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_55 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_54 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_53 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_52 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_51 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_50 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_49 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_48 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_47 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_46 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_45 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_44 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_43 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_42 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_41 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_40 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_39 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_38 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_37 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_36 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_35 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_34 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_33 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_32 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_31 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_30 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_28 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_27 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_26 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_25 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_24 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_23 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_22 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_21 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_20 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_19 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_18 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_17 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_15 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_14 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_13 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_12 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_11 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_10 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_9 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_8 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_7 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_6 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_5 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module CSTgen_CW4_NB32_7 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n3;

  pg_net_224 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_223 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_222 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_221 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_220 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_219 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_218 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_217 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_216 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_215 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_214 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_213 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_212 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_211 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_210 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_209 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_208 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_207 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_206 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_205 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_204 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_203 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_202 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_201 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_200 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_199 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_198 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_197 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_196 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_195 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_194 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_193 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_189 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_63 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_188 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_187 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_186 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_185 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_184 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_183 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_182 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_181 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_180 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_179 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_178 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_177 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_176 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_175 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_62 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_174 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_173 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_172 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_171 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_170 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_169 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_168 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_61 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_167 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_166 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_165 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_60 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_59 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_164 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_163 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_58 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_57 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_56 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_55 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(\matrixGen[0][0] ) );
endmodule


module CSTgen_CW4_NB32_6 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n3;

  pg_net_192 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_191 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_190 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_189 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_188 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_187 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_186 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_185 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_184 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_183 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_182 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_181 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_180 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_179 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_178 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_177 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_176 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_175 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_174 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_173 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_172 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_171 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_170 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_169 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_168 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_167 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_166 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_165 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_164 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_163 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_162 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_161 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_162 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_54 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_161 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_160 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_159 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_158 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_157 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_156 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_155 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_154 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_153 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_152 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_151 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_150 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_149 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_148 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_53 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_147 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_146 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_145 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_144 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_143 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_142 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_141 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_52 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_140 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_139 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_138 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_51 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_50 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_137 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_136 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_49 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_48 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_47 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_46 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(\matrixGen[0][0] ) );
endmodule


module CSTgen_CW4_NB32_5 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n3;

  pg_net_160 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_159 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_158 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_157 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_156 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_155 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_154 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_153 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_152 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_151 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_150 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_149 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_148 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_147 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_146 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_145 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_144 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_143 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_142 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_141 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_140 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_139 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_138 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_137 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_136 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_135 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_134 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_133 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_132 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_131 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_130 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_129 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_135 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_45 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_134 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_133 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_132 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_131 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_130 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_129 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_128 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_127 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_126 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_125 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_124 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_123 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_122 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_121 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_44 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_120 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_119 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_118 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_117 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_116 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_115 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_114 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_43 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_113 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_112 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_111 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_42 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_41 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_110 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_109 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_40 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_39 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_38 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_37 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(\matrixGen[0][0] ) );
endmodule


module CSTgen_CW4_NB32_3 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n3;

  pg_net_96 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_95 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_94 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_93 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_92 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_91 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_90 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_89 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_88 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_87 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_86 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_85 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_84 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_83 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_82 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_81 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_80 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_79 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_78 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_77 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_76 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_75 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_74 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_73 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_72 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_71 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_70 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_69 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_68 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_67 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_66 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_65 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_81 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_27 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_80 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_79 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_78 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_77 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_76 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_75 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_74 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_73 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_72 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_71 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_70 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_69 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_68 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_67 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_26 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_66 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_65 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_64 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_63 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_62 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_61 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_60 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_25 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_59 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_58 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_57 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_24 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_23 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_56 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_55 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_22 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_21 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_20 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_19 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(\matrixGen[0][0] ) );
endmodule


module MUX21_generic_NB32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109;

  INV_X1 U1 ( .A(n76), .ZN(n67) );
  BUF_X1 U2 ( .A(n77), .Z(n68) );
  BUF_X1 U3 ( .A(n77), .Z(n69) );
  BUF_X1 U4 ( .A(n68), .Z(n75) );
  BUF_X1 U5 ( .A(n73), .Z(n74) );
  BUF_X1 U6 ( .A(n77), .Z(n73) );
  BUF_X1 U7 ( .A(n77), .Z(n72) );
  BUF_X1 U8 ( .A(n74), .Z(n70) );
  BUF_X1 U9 ( .A(n77), .Z(n71) );
  BUF_X1 U10 ( .A(n77), .Z(n76) );
  INV_X1 U11 ( .A(SEL), .ZN(n77) );
  INV_X1 U12 ( .A(n104), .ZN(Y[4]) );
  AOI22_X1 U13 ( .A1(A[4]), .A2(SEL), .B1(B[4]), .B2(n69), .ZN(n104) );
  INV_X1 U14 ( .A(n106), .ZN(Y[6]) );
  AOI22_X1 U15 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(n68), .ZN(n106) );
  INV_X1 U16 ( .A(n108), .ZN(Y[8]) );
  AOI22_X1 U17 ( .A1(A[8]), .A2(SEL), .B1(B[8]), .B2(n68), .ZN(n108) );
  INV_X1 U18 ( .A(n103), .ZN(Y[3]) );
  AOI22_X1 U19 ( .A1(A[3]), .A2(SEL), .B1(B[3]), .B2(n69), .ZN(n103) );
  INV_X1 U20 ( .A(n105), .ZN(Y[5]) );
  AOI22_X1 U21 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(n69), .ZN(n105) );
  INV_X1 U22 ( .A(n107), .ZN(Y[7]) );
  AOI22_X1 U23 ( .A1(A[7]), .A2(SEL), .B1(B[7]), .B2(n68), .ZN(n107) );
  INV_X1 U24 ( .A(n102), .ZN(Y[31]) );
  AOI22_X1 U25 ( .A1(A[31]), .A2(SEL), .B1(B[31]), .B2(n69), .ZN(n102) );
  INV_X1 U26 ( .A(n101), .ZN(Y[30]) );
  AOI22_X1 U27 ( .A1(A[30]), .A2(n67), .B1(B[30]), .B2(n70), .ZN(n101) );
  AOI22_X1 U28 ( .A1(SEL), .A2(A[9]), .B1(B[9]), .B2(n68), .ZN(n109) );
  INV_X1 U29 ( .A(n91), .ZN(Y[21]) );
  AOI22_X1 U30 ( .A1(A[21]), .A2(n67), .B1(B[21]), .B2(n72), .ZN(n91) );
  INV_X1 U31 ( .A(n98), .ZN(Y[28]) );
  AOI22_X1 U32 ( .A1(A[28]), .A2(n67), .B1(B[28]), .B2(n70), .ZN(n98) );
  INV_X1 U33 ( .A(n90), .ZN(Y[20]) );
  AOI22_X1 U34 ( .A1(A[20]), .A2(n67), .B1(B[20]), .B2(n72), .ZN(n90) );
  INV_X1 U35 ( .A(n94), .ZN(Y[24]) );
  AOI22_X1 U36 ( .A1(A[24]), .A2(n67), .B1(B[24]), .B2(n71), .ZN(n94) );
  INV_X1 U37 ( .A(n95), .ZN(Y[25]) );
  AOI22_X1 U38 ( .A1(A[25]), .A2(n67), .B1(B[25]), .B2(n71), .ZN(n95) );
  INV_X1 U39 ( .A(n96), .ZN(Y[26]) );
  AOI22_X1 U40 ( .A1(A[26]), .A2(n67), .B1(B[26]), .B2(n71), .ZN(n96) );
  INV_X1 U41 ( .A(n97), .ZN(Y[27]) );
  AOI22_X1 U42 ( .A1(A[27]), .A2(n67), .B1(B[27]), .B2(n71), .ZN(n97) );
  INV_X1 U43 ( .A(n81), .ZN(Y[12]) );
  AOI22_X1 U44 ( .A1(A[12]), .A2(SEL), .B1(B[12]), .B2(n75), .ZN(n81) );
  INV_X1 U45 ( .A(n83), .ZN(Y[14]) );
  AOI22_X1 U46 ( .A1(A[14]), .A2(SEL), .B1(B[14]), .B2(n74), .ZN(n83) );
  INV_X1 U47 ( .A(n100), .ZN(Y[2]) );
  AOI22_X1 U48 ( .A1(A[2]), .A2(n67), .B1(B[2]), .B2(n70), .ZN(n100) );
  INV_X1 U49 ( .A(n89), .ZN(Y[1]) );
  AOI22_X1 U50 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n73), .ZN(n89) );
  INV_X1 U51 ( .A(n82), .ZN(Y[13]) );
  AOI22_X1 U52 ( .A1(A[13]), .A2(SEL), .B1(B[13]), .B2(n74), .ZN(n82) );
  INV_X1 U53 ( .A(n79), .ZN(Y[10]) );
  AOI22_X1 U54 ( .A1(A[10]), .A2(SEL), .B1(B[10]), .B2(n75), .ZN(n79) );
  INV_X1 U55 ( .A(n80), .ZN(Y[11]) );
  AOI22_X1 U56 ( .A1(A[11]), .A2(SEL), .B1(B[11]), .B2(n75), .ZN(n80) );
  INV_X1 U57 ( .A(n78), .ZN(Y[0]) );
  AOI22_X1 U58 ( .A1(A[0]), .A2(n67), .B1(B[0]), .B2(n75), .ZN(n78) );
  INV_X1 U59 ( .A(n87), .ZN(Y[18]) );
  AOI22_X1 U60 ( .A1(A[18]), .A2(SEL), .B1(B[18]), .B2(n73), .ZN(n87) );
  INV_X1 U61 ( .A(n92), .ZN(Y[22]) );
  AOI22_X1 U62 ( .A1(A[22]), .A2(n67), .B1(B[22]), .B2(n72), .ZN(n92) );
  INV_X1 U63 ( .A(n86), .ZN(Y[17]) );
  AOI22_X1 U64 ( .A1(A[17]), .A2(SEL), .B1(B[17]), .B2(n73), .ZN(n86) );
  INV_X1 U65 ( .A(n85), .ZN(Y[16]) );
  AOI22_X1 U66 ( .A1(A[16]), .A2(SEL), .B1(B[16]), .B2(n74), .ZN(n85) );
  INV_X1 U67 ( .A(n93), .ZN(Y[23]) );
  AOI22_X1 U68 ( .A1(A[23]), .A2(n67), .B1(B[23]), .B2(n72), .ZN(n93) );
  INV_X1 U69 ( .A(n84), .ZN(Y[15]) );
  AOI22_X1 U70 ( .A1(A[15]), .A2(SEL), .B1(B[15]), .B2(n74), .ZN(n84) );
  INV_X1 U71 ( .A(n88), .ZN(Y[19]) );
  AOI22_X1 U72 ( .A1(A[19]), .A2(SEL), .B1(B[19]), .B2(n73), .ZN(n88) );
  INV_X1 U73 ( .A(n99), .ZN(Y[29]) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n67), .B1(B[29]), .B2(n70), .ZN(n99) );
  INV_X1 U75 ( .A(n109), .ZN(Y[9]) );
endmodule


module FD_NB32_4 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n35, n69, n70, n71;
  assign n35 = RESET;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n71), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n71), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n71), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n71), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n71), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n71), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n71), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n71), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n69), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n69), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n69), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n69), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n69), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n69), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n69), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n69), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n69), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n69), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n69), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n69), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n70), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n70), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n70), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n70), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n70), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n70), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n70), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n70), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n70), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n70), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n70), .Q(Q[0]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n70), .Q(Q[9]) );
  BUF_X1 U3 ( .A(n35), .Z(n70) );
  BUF_X1 U4 ( .A(n35), .Z(n69) );
  BUF_X1 U5 ( .A(n35), .Z(n71) );
endmodule


module FD_NB32_3 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n35, n68, n69, n70;
  assign n35 = RESET;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n70), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n70), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n70), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n70), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n70), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n70), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n70), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n70), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n68), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n68), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n68), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n68), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n68), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n68), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n68), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n68), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n68), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n68), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n68), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n68), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n69), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n69), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n69), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n69), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n69), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n69), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n69), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n69), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n69), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n69), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n69), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n69), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n35), .Z(n69) );
  BUF_X1 U4 ( .A(n35), .Z(n68) );
  BUF_X1 U5 ( .A(n35), .Z(n70) );
endmodule


module FD_NB32_2 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n35, n68, n69, n70;
  assign n35 = RESET;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n70), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n70), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n70), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n70), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n70), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n70), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n70), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n70), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n68), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n68), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n68), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n68), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n68), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n68), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n68), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n68), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n68), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n68), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n68), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n68), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n69), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n69), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n69), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n69), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n69), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n69), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n69), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n69), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n69), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n69), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n69), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n69), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n35), .Z(n69) );
  BUF_X1 U4 ( .A(n35), .Z(n68) );
  BUF_X1 U5 ( .A(n35), .Z(n70) );
endmodule


module FD_NB32_1 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n35, n68, n69, n70;
  assign n35 = RESET;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n70), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n70), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n70), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n70), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n70), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n70), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n70), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n70), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n68), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n68), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n68), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n68), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n68), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n68), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n68), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n68), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n68), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n68), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n68), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n68), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n69), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n69), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n69), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n69), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n69), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n69), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n69), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n69), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n69), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n69), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n69), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n69), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n35), .Z(n69) );
  BUF_X1 U4 ( .A(n35), .Z(n68) );
  BUF_X1 U5 ( .A(n35), .Z(n70) );
endmodule


module FD_INJ_NB32_1 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n38, n71, n72, n73, n74, n75, n76;
  wire   [31:0] TMP_D;
  assign n38 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n76), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n76), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n76), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n76), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n76), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n76), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n76), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n76), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n74), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n74), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n74), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n74), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n74), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n74), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n74), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n74), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n74), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n74), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n74), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n74), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n75), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n75), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n75), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n75), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n75), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n75), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n75), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n75), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n75), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n75), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n75), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n75), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n38), .Z(n75) );
  BUF_X1 U4 ( .A(n38), .Z(n74) );
  BUF_X1 U5 ( .A(n38), .Z(n76) );
  BUF_X1 U6 ( .A(INJ_ZERO), .Z(n71) );
  BUF_X1 U7 ( .A(INJ_ZERO), .Z(n72) );
  BUF_X1 U8 ( .A(INJ_ZERO), .Z(n73) );
  AND2_X1 U9 ( .A1(D[0]), .A2(n71), .ZN(TMP_D[0]) );
  AND2_X1 U10 ( .A1(D[1]), .A2(n71), .ZN(TMP_D[1]) );
  AND2_X1 U11 ( .A1(D[2]), .A2(n72), .ZN(TMP_D[2]) );
  AND2_X1 U12 ( .A1(D[10]), .A2(n71), .ZN(TMP_D[10]) );
  AND2_X1 U13 ( .A1(D[11]), .A2(n71), .ZN(TMP_D[11]) );
  AND2_X1 U14 ( .A1(D[12]), .A2(n71), .ZN(TMP_D[12]) );
  AND2_X1 U15 ( .A1(D[13]), .A2(n71), .ZN(TMP_D[13]) );
  AND2_X1 U16 ( .A1(D[14]), .A2(n71), .ZN(TMP_D[14]) );
  AND2_X1 U17 ( .A1(D[15]), .A2(n71), .ZN(TMP_D[15]) );
  AND2_X1 U18 ( .A1(D[16]), .A2(n71), .ZN(TMP_D[16]) );
  AND2_X1 U19 ( .A1(D[17]), .A2(n71), .ZN(TMP_D[17]) );
  AND2_X1 U20 ( .A1(D[18]), .A2(n71), .ZN(TMP_D[18]) );
  AND2_X1 U21 ( .A1(D[19]), .A2(n71), .ZN(TMP_D[19]) );
  AND2_X1 U22 ( .A1(D[20]), .A2(n72), .ZN(TMP_D[20]) );
  AND2_X1 U23 ( .A1(D[21]), .A2(n72), .ZN(TMP_D[21]) );
  AND2_X1 U24 ( .A1(D[22]), .A2(n72), .ZN(TMP_D[22]) );
  AND2_X1 U25 ( .A1(D[23]), .A2(n72), .ZN(TMP_D[23]) );
  AND2_X1 U26 ( .A1(D[24]), .A2(n72), .ZN(TMP_D[24]) );
  AND2_X1 U27 ( .A1(D[25]), .A2(n72), .ZN(TMP_D[25]) );
  AND2_X1 U28 ( .A1(D[26]), .A2(n72), .ZN(TMP_D[26]) );
  AND2_X1 U29 ( .A1(D[27]), .A2(n72), .ZN(TMP_D[27]) );
  AND2_X1 U30 ( .A1(D[28]), .A2(n72), .ZN(TMP_D[28]) );
  AND2_X1 U31 ( .A1(D[29]), .A2(n72), .ZN(TMP_D[29]) );
  AND2_X1 U32 ( .A1(D[30]), .A2(n72), .ZN(TMP_D[30]) );
  AND2_X1 U33 ( .A1(n73), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U34 ( .A1(D[3]), .A2(n73), .ZN(TMP_D[3]) );
  AND2_X1 U35 ( .A1(D[4]), .A2(n73), .ZN(TMP_D[4]) );
  AND2_X1 U36 ( .A1(D[5]), .A2(n73), .ZN(TMP_D[5]) );
  AND2_X1 U37 ( .A1(D[6]), .A2(n73), .ZN(TMP_D[6]) );
  AND2_X1 U38 ( .A1(D[7]), .A2(n73), .ZN(TMP_D[7]) );
  AND2_X1 U39 ( .A1(D[8]), .A2(n73), .ZN(TMP_D[8]) );
  AND2_X1 U40 ( .A1(D[31]), .A2(n73), .ZN(TMP_D[31]) );
endmodule


module FD_INJ_NB1_2 ( CK, RESET, INJ_ZERO, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   \TMP_D[0] ;

  DFFR_X1 \Q_reg[0]  ( .D(\TMP_D[0] ), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[0]), .ZN(\TMP_D[0] ) );
endmodule


module FD_INJ_NB1_1 ( CK, RESET, INJ_ZERO, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   \TMP_D[0] ;

  DFFR_X1 \Q_reg[0]  ( .D(\TMP_D[0] ), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[0]), .ZN(\TMP_D[0] ) );
endmodule


module FD_NB4_1 ( CK, RESET, D, Q );
  input [3:0] D;
  output [3:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB3_1 ( CK, RESET, D, Q );
  input [2:0] D;
  output [2:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB2_3 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB2_2 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB2_1 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_22 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_21 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_20 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_19 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_18 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_17 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_16 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_15 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X2 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_14 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_13 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_12 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_11 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_10 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_9 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_8 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_7 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_6 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_5 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_4 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_3 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_2 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_1 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB11_1 ( CK, RESET, D, Q );
  input [10:0] D;
  output [10:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(RESET), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(RESET), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(RESET), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(RESET), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(RESET), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_3 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_2 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_1 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module carry_sel_bk_NB4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  OAI22_X1 U3 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U4 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  INV_X1 U5 ( .A(B[1]), .ZN(n18) );
  NAND2_X1 U6 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U7 ( .A(n21), .ZN(n26) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  AOI22_X1 U10 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U13 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U14 ( .A(A[1]), .ZN(n17) );
  OR2_X1 U15 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  OAI22_X1 U16 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  OAI22_X1 U17 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  OAI22_X1 U18 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
endmodule


module carry_sel_bk_NB4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  OAI22_X1 U3 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U4 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  INV_X1 U5 ( .A(B[1]), .ZN(n18) );
  NAND2_X1 U6 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U7 ( .A(n21), .ZN(n26) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  AOI22_X1 U10 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U13 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U14 ( .A(A[1]), .ZN(n17) );
  OR2_X1 U15 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  OAI22_X1 U16 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U17 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  OAI22_X1 U18 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
endmodule


module carry_sel_bk_NB4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NOR2_X1 U7 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  NOR2_X1 U9 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  INV_X1 U10 ( .A(B[1]), .ZN(n18) );
  AOI22_X1 U11 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  AOI22_X1 U12 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  XNOR2_X1 U13 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OR2_X1 U14 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  OAI22_X1 U15 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  OAI22_X1 U16 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  OAI22_X1 U17 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  OAI22_X1 U3 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U4 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  INV_X1 U5 ( .A(B[1]), .ZN(n18) );
  NAND2_X1 U6 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U7 ( .A(n21), .ZN(n26) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  AOI22_X1 U10 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  AOI22_X1 U11 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U13 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OR2_X1 U14 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  OAI22_X1 U15 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U16 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  OAI22_X1 U17 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n46, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n46), .B(n25), .Z(S[0]) );
  OAI22_X1 U2 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U3 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  INV_X1 U4 ( .A(B[1]), .ZN(n18) );
  NAND2_X1 U5 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U6 ( .A(n21), .ZN(n26) );
  NOR2_X1 U7 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  AOI22_X1 U10 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U11 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U12 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OR2_X1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  OAI22_X1 U14 ( .A1(n46), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U15 ( .A1(n46), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  OAI22_X1 U16 ( .A1(n46), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  INV_X1 U17 ( .A(Ci), .ZN(n46) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_13 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  INV_X1 U7 ( .A(B[1]), .ZN(n18) );
  OAI22_X1 U8 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U10 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U17 ( .A(A[1]), .ZN(n17) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
endmodule


module carry_sel_bk_NB4_16 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n46, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n46), .B(n25), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U3 ( .A(n21), .ZN(n26) );
  OAI22_X1 U4 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U6 ( .A1(n46), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U7 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U8 ( .A1(n46), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U9 ( .A1(n46), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U10 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U11 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  AOI22_X1 U12 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U14 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U15 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U17 ( .A(Ci), .ZN(n46) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_18 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U6 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U7 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U8 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  OAI22_X1 U9 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U10 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  AOI22_X1 U11 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U12 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  OAI22_X1 U14 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  NOR2_X1 U15 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U16 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U17 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U18 ( .A(A[1]), .ZN(n17) );
endmodule


module carry_sel_bk_NB4_22 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U7 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NAND2_X1 U9 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  NOR2_X1 U10 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  INV_X1 U11 ( .A(B[1]), .ZN(n18) );
  OAI22_X1 U12 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U13 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U15 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_24 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n46, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n46), .B(n25), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U3 ( .A(n21), .ZN(n26) );
  OAI22_X1 U4 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U6 ( .A1(n46), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U7 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U8 ( .A1(n46), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U9 ( .A1(n46), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U10 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U11 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NAND2_X1 U12 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U15 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U17 ( .A(Ci), .ZN(n46) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_30 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  INV_X1 U7 ( .A(B[1]), .ZN(n18) );
  OAI22_X1 U8 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U10 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U17 ( .A(A[1]), .ZN(n17) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
endmodule


module blockPG_104 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module carry_sel_bk_NB4_35 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U6 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U7 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U8 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  OAI22_X1 U9 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U10 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  AOI22_X1 U11 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U12 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  OAI22_X1 U14 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  NOR2_X1 U15 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U16 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U17 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U18 ( .A(A[1]), .ZN(n17) );
endmodule


module carry_sel_bk_NB4_39 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U7 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  NOR2_X1 U8 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U9 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U10 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U11 ( .A(B[1]), .ZN(n18) );
  OAI22_X1 U12 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U13 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U15 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_40 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n46, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n46), .B(n25), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U3 ( .A(n21), .ZN(n26) );
  OAI22_X1 U4 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U6 ( .A1(n46), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U7 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U8 ( .A1(n46), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U9 ( .A1(n46), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U10 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U11 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  AOI22_X1 U12 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND2_X1 U14 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U15 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U17 ( .A(Ci), .ZN(n46) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_41 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  NOR2_X1 U5 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U7 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OAI22_X1 U9 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U10 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U11 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U12 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U16 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_42 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  NOR2_X1 U5 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U7 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OAI22_X1 U9 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U10 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U11 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U12 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U16 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_43 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U3 ( .A(n21), .ZN(n26) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NOR2_X1 U5 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U7 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OAI22_X1 U9 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U10 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U11 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U12 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U16 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_47 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U7 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U9 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U12 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U13 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U16 ( .A(A[1]), .ZN(n17) );
  INV_X1 U17 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
endmodule


module carry_sel_bk_NB4_48 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n48, n49;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n48), .B(n25), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U3 ( .A(n21), .ZN(n26) );
  OAI22_X1 U4 ( .A1(n49), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U5 ( .A1(n49), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U6 ( .A1(n48), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U7 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U8 ( .A1(n48), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U9 ( .A1(n48), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U10 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U11 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NAND2_X1 U14 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U15 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U17 ( .A(Ci), .ZN(n48) );
  INV_X1 U18 ( .A(A[1]), .ZN(n49) );
endmodule


module carry_sel_bk_NB4_50 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NOR2_X1 U7 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OAI22_X1 U9 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U10 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U11 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U12 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U16 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_51 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NOR2_X1 U7 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OAI22_X1 U9 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U10 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U11 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U12 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U13 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U16 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_52 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  NOR2_X1 U5 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  OAI22_X1 U6 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U7 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U9 ( .A(A[1]), .ZN(n17) );
  OAI22_X1 U10 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U12 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U13 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U14 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NOR2_X1 U16 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  INV_X1 U17 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
endmodule


module carry_sel_bk_NB4_56 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U3 ( .A(n21), .ZN(n26) );
  OAI22_X1 U4 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U5 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  NOR2_X1 U6 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  INV_X1 U7 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U8 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  INV_X1 U9 ( .A(A[1]), .ZN(n17) );
  OAI22_X1 U10 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U11 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U12 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U13 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U14 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U15 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U16 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  INV_X1 U17 ( .A(B[1]), .ZN(n18) );
  OR2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
endmodule


module carry_sel_bk_NB4_59 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U7 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U9 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NOR2_X1 U14 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U17 ( .A(B[1]), .ZN(n18) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_60 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n47;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n47), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n47), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U7 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U8 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U9 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U10 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U11 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NOR2_X1 U14 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NAND2_X1 U15 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OR2_X1 U16 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U17 ( .A(B[1]), .ZN(n18) );
  INV_X1 U18 ( .A(A[1]), .ZN(n47) );
endmodule


module carry_sel_bk_NB4_62 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  INV_X1 U3 ( .A(A[1]), .ZN(n17) );
  NAND2_X1 U4 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U5 ( .A(n21), .ZN(n26) );
  OAI22_X1 U6 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U7 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U8 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U10 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(B[1]), .ZN(n18) );
endmodule


module carry_sel_bk_NB4_63 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(Ci), .ZN(n5) );
  INV_X1 U3 ( .A(A[1]), .ZN(n17) );
  NAND2_X1 U4 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U5 ( .A(n21), .ZN(n26) );
  OAI22_X1 U6 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U7 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  OAI22_X1 U8 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U10 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(B[1]), .ZN(n18) );
endmodule


module carry_sel_bk_NB4_64 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26;

  XOR2_X1 U19 ( .A(n8), .B(n9), .Z(n7) );
  XOR2_X1 U20 ( .A(n12), .B(n9), .Z(n6) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U22 ( .A(n10), .B(n16), .Z(n15) );
  XOR2_X1 U23 ( .A(n13), .B(n16), .Z(n14) );
  XOR2_X1 U24 ( .A(n20), .B(n24), .Z(n23) );
  XOR2_X1 U25 ( .A(n21), .B(n24), .Z(n22) );
  XOR2_X1 U26 ( .A(A[1]), .B(B[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(n5), .B(n25), .Z(S[0]) );
  INV_X1 U2 ( .A(A[1]), .ZN(n17) );
  NAND2_X1 U3 ( .A1(n26), .A2(n20), .ZN(n25) );
  INV_X1 U4 ( .A(n21), .ZN(n26) );
  OAI22_X1 U5 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n10) );
  OAI22_X1 U6 ( .A1(n17), .A2(n18), .B1(n21), .B2(n19), .ZN(n13) );
  INV_X1 U7 ( .A(Ci), .ZN(n5) );
  OAI22_X1 U8 ( .A1(n5), .A2(n14), .B1(Ci), .B2(n15), .ZN(S[2]) );
  XNOR2_X1 U9 ( .A(A[2]), .B(B[2]), .ZN(n16) );
  OAI22_X1 U10 ( .A1(n5), .A2(n22), .B1(Ci), .B2(n23), .ZN(S[1]) );
  OAI22_X1 U11 ( .A1(n5), .A2(n6), .B1(Ci), .B2(n7), .ZN(S[3]) );
  AOI22_X1 U12 ( .A1(n10), .A2(n11), .B1(B[2]), .B2(A[2]), .ZN(n8) );
  NOR2_X1 U13 ( .A1(A[0]), .A2(B[0]), .ZN(n21) );
  NOR2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(B[2]), .B1(n13), .B2(n11), .ZN(n12) );
  NAND2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n20) );
  OR2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  INV_X1 U18 ( .A(B[1]), .ZN(n18) );
endmodule


module blockPG_201 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
endmodule


module sum_gen_Nrca4_NB32_1 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_8 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  carry_sel_bk_NB4_7 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  carry_sel_bk_NB4_6 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  carry_sel_bk_NB4_5 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_4 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_3 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_2 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_1 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_1 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n2;

  pg_net_32 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_31 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_30 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_29 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_28 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_27 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_26 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_25 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_24 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_23 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_22 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_21 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_20 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_19 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_18 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_17 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_16 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_15 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_14 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_13 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_12 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_11 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_10 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_9 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_8 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_7 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_6 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_5 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_4 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_3 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_2 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_1 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_27 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_9 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_26 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_25 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_24 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_23 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_22 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_21 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_20 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_19 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_18 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_17 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_16 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_15 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_14 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_13 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_8 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_12 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_11 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_10 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_9 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_8 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_7 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_6 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_7 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_5 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_4 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_3 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_6 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_5 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_2 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_1 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_4 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_3 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_2 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_1 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(\matrixGen[0][0] ) );
endmodule


module sum_gen_Nrca4_NB32_2 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_16 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_15 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_14 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_13 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_12 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_11 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_10 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_9 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_2 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n2;

  pg_net_64 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_63 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_62 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_61 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_60 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_59 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_58 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_57 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_56 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_55 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_54 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_53 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_52 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_51 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_50 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_49 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_48 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_47 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_46 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_45 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_44 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_43 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_42 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_41 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_40 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_39 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_38 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_37 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_36 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_35 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_34 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_33 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_54 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_18 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_53 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_52 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_51 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_50 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_49 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_48 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_47 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_46 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_45 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_44 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_43 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_42 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_41 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_40 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_17 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_39 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_38 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_37 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_36 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_35 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_34 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_33 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_16 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_32 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_31 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_30 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_15 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_14 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_29 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_28 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_13 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_12 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_11 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_10 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(\matrixGen[0][0] ) );
endmodule


module sum_gen_Nrca4_NB32_3 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_24 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_23 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_22 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_21 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_20 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_19 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_18 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_17 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_4 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_32 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_31 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_30 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_29 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_28 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_27 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_26 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_25 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_4 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n2;

  pg_net_128 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_127 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_126 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_125 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_124 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_123 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_122 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_121 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_120 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_119 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_118 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_117 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_116 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_115 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_114 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_113 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_112 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_111 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_110 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_109 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_108 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_107 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_106 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_105 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_104 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_103 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_102 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_101 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_100 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_99 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_98 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_97 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_108 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_36 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_107 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_106 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_105 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_104 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_103 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_102 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_101 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_100 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_99 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_98 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_97 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_96 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_95 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_94 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_35 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_93 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_92 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_91 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_90 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_89 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_88 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_87 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_34 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_86 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), 
        .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_85 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), 
        .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_84 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), 
        .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_33 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_32 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_83 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_82 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), 
        .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_31 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_30 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_29 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_28 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(\matrixGen[0][0] ) );
endmodule


module sum_gen_Nrca4_NB32_5 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_40 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_39 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_38 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_37 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_36 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_35 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_34 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_33 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_6 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_48 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_47 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_46 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_45 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_44 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_43 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_42 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_41 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_7 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_56 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_55 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_54 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_53 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_52 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_51 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_50 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_49 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sum_gen_Nrca4_NB32_8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_64 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  carry_sel_bk_NB4_63 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_62 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_61 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_60 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_59 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_58 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_57 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_8 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[0][0] , \matrixGen[1][31] , \matrixGen[1][29] ,
         \matrixGen[1][27] , \matrixGen[1][25] , \matrixGen[1][23] ,
         \matrixGen[1][21] , \matrixGen[1][19] , \matrixGen[1][17] ,
         \matrixGen[1][15] , \matrixGen[1][13] , \matrixGen[1][11] ,
         \matrixGen[1][9] , \matrixGen[1][7] , \matrixGen[1][5] ,
         \matrixGen[1][3] , \matrixGen[1][1] , \matrixGen[2][31] ,
         \matrixGen[2][27] , \matrixGen[2][23] , \matrixGen[2][19] ,
         \matrixGen[2][15] , \matrixGen[2][11] , \matrixGen[2][7] ,
         \matrixGen[3][31] , \matrixGen[3][23] , \matrixGen[3][15] ,
         \matrixGen[4][31] , \matrixGen[4][27] , n2;

  pg_net_256 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp)
         );
  pg_net_255 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_254 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_253 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_252 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_251 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_250 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_249 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_248 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_247 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_246 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_245 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_244 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_243 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_242 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_241 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_240 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_239 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_238 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_237 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_236 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_235 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_234 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_233 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_232 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_231 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_230 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_229 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_228 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_227 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_226 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_225 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_216 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_72 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(\matrixGen[0][0] ), .Pik(
        \matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_215 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_214 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_213 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_212 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_211 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_210 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_209 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_208 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_207 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_206 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_205 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_204 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_203 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_202 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_71 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(C[0]) );
  blockPG_201 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_200 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_199 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_198 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_197 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_196 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_195 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_70 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(C[0]), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_194 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_193 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_192 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_69 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_68 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_191 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_190 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_67 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_66 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_65 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_64 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  AOI21_X1 U1 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(\matrixGen[0][0] ) );
endmodule


module carry_sel_bk_NB4_65 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31;

  XOR2_X1 U29 ( .A(n18), .B(n19), .Z(S[2]) );
  XOR2_X1 U30 ( .A(n9), .B(n30), .Z(S[0]) );
  OAI22_X2 U2 ( .A1(n24), .A2(n25), .B1(n26), .B2(n27), .ZN(S[1]) );
  NAND2_X1 U3 ( .A1(n31), .A2(n23), .ZN(n30) );
  INV_X1 U4 ( .A(n21), .ZN(n31) );
  INV_X1 U5 ( .A(n27), .ZN(n24) );
  NAND2_X1 U6 ( .A1(n29), .A2(n22), .ZN(n27) );
  OAI21_X1 U7 ( .B1(n20), .B2(n23), .A(n22), .ZN(n15) );
  OAI21_X1 U8 ( .B1(n20), .B2(n21), .A(n22), .ZN(n13) );
  INV_X1 U9 ( .A(n20), .ZN(n29) );
  XNOR2_X1 U10 ( .A(n10), .B(n11), .ZN(n8) );
  XNOR2_X1 U11 ( .A(n14), .B(n10), .ZN(n7) );
  XNOR2_X1 U12 ( .A(B[3]), .B(A[3]), .ZN(n10) );
  XNOR2_X1 U13 ( .A(B[2]), .B(A[2]), .ZN(n19) );
  OAI22_X1 U14 ( .A1(n12), .A2(B[2]), .B1(n13), .B2(A[2]), .ZN(n11) );
  AND2_X1 U15 ( .A1(A[2]), .A2(n13), .ZN(n12) );
  NOR2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  NOR2_X1 U17 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  NAND2_X1 U18 ( .A1(B[0]), .A2(A[0]), .ZN(n23) );
  NAND2_X1 U19 ( .A1(B[1]), .A2(A[1]), .ZN(n22) );
  AOI21_X1 U20 ( .B1(n15), .B2(A[2]), .A(n16), .ZN(n14) );
  INV_X1 U21 ( .A(n17), .ZN(n16) );
  OAI21_X1 U22 ( .B1(A[2]), .B2(n15), .A(B[2]), .ZN(n17) );
  OAI21_X1 U23 ( .B1(Ci), .B2(n15), .A(n13), .ZN(n18) );
  OAI22_X1 U24 ( .A1(Ci), .A2(n7), .B1(n8), .B2(n9), .ZN(S[3]) );
  INV_X1 U25 ( .A(n28), .ZN(n25) );
  AOI21_X1 U26 ( .B1(n23), .B2(n9), .A(n21), .ZN(n26) );
  INV_X1 U27 ( .A(Ci), .ZN(n9) );
  OAI21_X1 U28 ( .B1(n9), .B2(n21), .A(n23), .ZN(n28) );
endmodule


module carry_sel_bk_NB4_66 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29;

  XOR2_X1 U28 ( .A(n16), .B(n17), .Z(S[2]) );
  XOR2_X1 U29 ( .A(n8), .B(n28), .Z(S[0]) );
  OAI22_X2 U2 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(S[1]) );
  NAND2_X1 U3 ( .A1(n29), .A2(n21), .ZN(n28) );
  INV_X1 U4 ( .A(n19), .ZN(n29) );
  INV_X1 U5 ( .A(n25), .ZN(n22) );
  NAND2_X1 U6 ( .A1(n27), .A2(n20), .ZN(n25) );
  OAI21_X1 U7 ( .B1(n18), .B2(n21), .A(n20), .ZN(n15) );
  OAI21_X1 U8 ( .B1(n18), .B2(n19), .A(n20), .ZN(n11) );
  OAI21_X1 U9 ( .B1(n11), .B2(n12), .A(n13), .ZN(n10) );
  OAI21_X1 U10 ( .B1(n12), .B2(n15), .A(n13), .ZN(n14) );
  INV_X1 U11 ( .A(n18), .ZN(n27) );
  XNOR2_X1 U12 ( .A(n9), .B(n10), .ZN(n7) );
  XNOR2_X1 U13 ( .A(n14), .B(n9), .ZN(n6) );
  XNOR2_X1 U14 ( .A(B[3]), .B(A[3]), .ZN(n9) );
  XNOR2_X1 U15 ( .A(A[2]), .B(B[2]), .ZN(n17) );
  NOR2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n19) );
  NOR2_X1 U17 ( .A1(B[1]), .A2(A[1]), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  NAND2_X1 U19 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  AND2_X1 U20 ( .A1(B[2]), .A2(A[2]), .ZN(n12) );
  OR2_X1 U21 ( .A1(A[2]), .A2(B[2]), .ZN(n13) );
  OAI21_X1 U22 ( .B1(Ci), .B2(n15), .A(n11), .ZN(n16) );
  OAI22_X1 U23 ( .A1(Ci), .A2(n6), .B1(n7), .B2(n8), .ZN(S[3]) );
  AOI21_X1 U24 ( .B1(n21), .B2(n8), .A(n19), .ZN(n24) );
  OAI21_X1 U25 ( .B1(n8), .B2(n19), .A(n21), .ZN(n26) );
  INV_X1 U26 ( .A(Ci), .ZN(n8) );
  INV_X1 U27 ( .A(n26), .ZN(n23) );
endmodule


module carry_sel_bk_NB4_67 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n29, n30;

  XOR2_X1 U2 ( .A(Ci), .B(n30), .Z(S[0]) );
  AND2_X1 U3 ( .A1(n29), .A2(n21), .ZN(n30) );
  INV_X1 U4 ( .A(n19), .ZN(n29) );
  INV_X1 U5 ( .A(n25), .ZN(n22) );
  NAND2_X1 U6 ( .A1(n27), .A2(n20), .ZN(n25) );
  OAI21_X1 U7 ( .B1(n18), .B2(n21), .A(n20), .ZN(n15) );
  OAI21_X1 U8 ( .B1(n18), .B2(n19), .A(n20), .ZN(n11) );
  OAI21_X1 U9 ( .B1(n11), .B2(n12), .A(n13), .ZN(n10) );
  OAI21_X1 U10 ( .B1(n12), .B2(n15), .A(n13), .ZN(n14) );
  INV_X1 U11 ( .A(n18), .ZN(n27) );
  XNOR2_X1 U12 ( .A(n14), .B(n9), .ZN(n6) );
  XNOR2_X1 U13 ( .A(n9), .B(n10), .ZN(n7) );
  XNOR2_X1 U14 ( .A(B[3]), .B(A[3]), .ZN(n9) );
  XNOR2_X1 U15 ( .A(A[2]), .B(B[2]), .ZN(n17) );
  NOR2_X1 U16 ( .A1(B[0]), .A2(A[0]), .ZN(n19) );
  NOR2_X1 U17 ( .A1(B[1]), .A2(A[1]), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  NAND2_X1 U19 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  AND2_X1 U20 ( .A1(B[2]), .A2(A[2]), .ZN(n12) );
  OR2_X1 U21 ( .A1(A[2]), .A2(B[2]), .ZN(n13) );
  XOR2_X1 U22 ( .A(n16), .B(n17), .Z(S[2]) );
  OAI22_X1 U23 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(S[1]) );
  OAI21_X1 U24 ( .B1(Ci), .B2(n15), .A(n11), .ZN(n16) );
  INV_X1 U25 ( .A(Ci), .ZN(n8) );
  OAI22_X1 U26 ( .A1(n6), .A2(Ci), .B1(n7), .B2(n8), .ZN(S[3]) );
  INV_X1 U27 ( .A(n26), .ZN(n23) );
  AOI21_X1 U28 ( .B1(n21), .B2(n8), .A(n19), .ZN(n24) );
  OAI21_X1 U29 ( .B1(n8), .B2(n19), .A(n21), .ZN(n26) );
endmodule


module carry_sel_bk_NB4_68 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29;

  XOR2_X1 U28 ( .A(n16), .B(n17), .Z(S[2]) );
  XOR2_X1 U29 ( .A(n8), .B(n28), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n29), .A2(n21), .ZN(n28) );
  INV_X1 U3 ( .A(n19), .ZN(n29) );
  OAI22_X1 U4 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(S[1]) );
  INV_X1 U5 ( .A(n25), .ZN(n22) );
  NAND2_X1 U6 ( .A1(n27), .A2(n20), .ZN(n25) );
  OAI21_X1 U7 ( .B1(n18), .B2(n21), .A(n20), .ZN(n15) );
  OAI21_X1 U8 ( .B1(n18), .B2(n19), .A(n20), .ZN(n11) );
  OAI21_X1 U9 ( .B1(n11), .B2(n12), .A(n13), .ZN(n10) );
  OAI21_X1 U10 ( .B1(n12), .B2(n15), .A(n13), .ZN(n14) );
  INV_X1 U11 ( .A(n18), .ZN(n27) );
  INV_X1 U12 ( .A(n26), .ZN(n23) );
  XNOR2_X1 U13 ( .A(n9), .B(n10), .ZN(n7) );
  XNOR2_X1 U14 ( .A(n14), .B(n9), .ZN(n6) );
  XNOR2_X1 U15 ( .A(B[3]), .B(A[3]), .ZN(n9) );
  XNOR2_X1 U16 ( .A(A[2]), .B(B[2]), .ZN(n17) );
  NOR2_X1 U17 ( .A1(B[0]), .A2(A[0]), .ZN(n19) );
  NOR2_X1 U18 ( .A1(B[1]), .A2(A[1]), .ZN(n18) );
  NAND2_X1 U19 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  NAND2_X1 U20 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  AND2_X1 U21 ( .A1(B[2]), .A2(A[2]), .ZN(n12) );
  OR2_X1 U22 ( .A1(A[2]), .A2(B[2]), .ZN(n13) );
  AOI21_X1 U23 ( .B1(n21), .B2(n8), .A(n19), .ZN(n24) );
  OAI21_X1 U24 ( .B1(n8), .B2(n19), .A(n21), .ZN(n26) );
  OAI22_X1 U25 ( .A1(Ci), .A2(n6), .B1(n7), .B2(n8), .ZN(S[3]) );
  OAI21_X1 U26 ( .B1(Ci), .B2(n15), .A(n11), .ZN(n16) );
  INV_X1 U27 ( .A(Ci), .ZN(n8) );
endmodule


module carry_sel_bk_NB4_69 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31;

  XOR2_X1 U29 ( .A(n18), .B(n19), .Z(S[2]) );
  XOR2_X1 U30 ( .A(n8), .B(n30), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n17), .A2(n12), .ZN(n18) );
  NAND2_X1 U3 ( .A1(n31), .A2(n23), .ZN(n30) );
  INV_X1 U4 ( .A(n21), .ZN(n31) );
  OAI22_X1 U5 ( .A1(n24), .A2(n25), .B1(n26), .B2(n27), .ZN(S[1]) );
  INV_X1 U6 ( .A(n27), .ZN(n24) );
  NAND2_X1 U7 ( .A1(n29), .A2(n22), .ZN(n27) );
  OAI21_X1 U8 ( .B1(n20), .B2(n21), .A(n22), .ZN(n13) );
  AOI21_X1 U9 ( .B1(n16), .B2(n12), .A(n14), .ZN(n15) );
  AOI21_X1 U10 ( .B1(n12), .B2(n13), .A(n14), .ZN(n10) );
  OAI21_X1 U11 ( .B1(n20), .B2(n23), .A(n22), .ZN(n16) );
  INV_X1 U12 ( .A(n17), .ZN(n14) );
  INV_X1 U13 ( .A(n20), .ZN(n29) );
  XNOR2_X1 U14 ( .A(n15), .B(n11), .ZN(n7) );
  XNOR2_X1 U15 ( .A(n10), .B(n11), .ZN(n9) );
  XNOR2_X1 U16 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  NOR2_X1 U17 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  NAND2_X1 U18 ( .A1(B[0]), .A2(A[0]), .ZN(n23) );
  NAND2_X1 U19 ( .A1(B[2]), .A2(A[2]), .ZN(n17) );
  OR2_X1 U20 ( .A1(A[2]), .A2(B[2]), .ZN(n12) );
  NAND2_X1 U21 ( .A1(B[1]), .A2(A[1]), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  OAI21_X1 U23 ( .B1(Ci), .B2(n16), .A(n13), .ZN(n19) );
  INV_X1 U24 ( .A(Ci), .ZN(n8) );
  OAI22_X1 U25 ( .A1(Ci), .A2(n7), .B1(n8), .B2(n9), .ZN(S[3]) );
  INV_X1 U26 ( .A(n28), .ZN(n25) );
  AOI21_X1 U27 ( .B1(n23), .B2(n8), .A(n21), .ZN(n26) );
  OAI21_X1 U28 ( .B1(n8), .B2(n21), .A(n23), .ZN(n28) );
endmodule


module carry_sel_bk_NB4_70 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29;

  XOR2_X1 U28 ( .A(n16), .B(n17), .Z(S[2]) );
  XOR2_X1 U29 ( .A(n8), .B(n28), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n29), .A2(n21), .ZN(n28) );
  INV_X1 U3 ( .A(n19), .ZN(n29) );
  OAI22_X1 U4 ( .A1(n22), .A2(n23), .B1(n24), .B2(n25), .ZN(S[1]) );
  INV_X1 U5 ( .A(n25), .ZN(n22) );
  NAND2_X1 U6 ( .A1(n27), .A2(n20), .ZN(n25) );
  AOI21_X1 U7 ( .B1(n21), .B2(n8), .A(n19), .ZN(n24) );
  OAI21_X1 U8 ( .B1(n18), .B2(n21), .A(n20), .ZN(n15) );
  OAI21_X1 U9 ( .B1(n18), .B2(n19), .A(n20), .ZN(n11) );
  OAI21_X1 U10 ( .B1(n11), .B2(n12), .A(n13), .ZN(n10) );
  OAI21_X1 U11 ( .B1(n12), .B2(n15), .A(n13), .ZN(n14) );
  INV_X1 U12 ( .A(n18), .ZN(n27) );
  INV_X1 U13 ( .A(n26), .ZN(n23) );
  OAI21_X1 U14 ( .B1(n8), .B2(n19), .A(n21), .ZN(n26) );
  XNOR2_X1 U15 ( .A(n9), .B(n10), .ZN(n7) );
  XNOR2_X1 U16 ( .A(n14), .B(n9), .ZN(n6) );
  XNOR2_X1 U17 ( .A(B[3]), .B(A[3]), .ZN(n9) );
  NOR2_X1 U18 ( .A1(B[0]), .A2(A[0]), .ZN(n19) );
  NAND2_X1 U19 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  OR2_X1 U20 ( .A1(A[2]), .A2(B[2]), .ZN(n13) );
  AND2_X1 U21 ( .A1(B[2]), .A2(A[2]), .ZN(n12) );
  XNOR2_X1 U22 ( .A(A[2]), .B(B[2]), .ZN(n17) );
  OAI22_X1 U23 ( .A1(Ci), .A2(n6), .B1(n7), .B2(n8), .ZN(S[3]) );
  OAI21_X1 U24 ( .B1(Ci), .B2(n15), .A(n11), .ZN(n16) );
  INV_X1 U25 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  NOR2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n18) );
endmodule


module carry_sel_bk_NB4_71 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31;

  XOR2_X1 U29 ( .A(n18), .B(n19), .Z(S[2]) );
  XOR2_X1 U30 ( .A(n8), .B(n30), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n17), .A2(n12), .ZN(n18) );
  NAND2_X1 U3 ( .A1(n31), .A2(n23), .ZN(n30) );
  INV_X1 U4 ( .A(n21), .ZN(n31) );
  OAI22_X1 U5 ( .A1(n24), .A2(n25), .B1(n26), .B2(n27), .ZN(S[1]) );
  INV_X1 U6 ( .A(n27), .ZN(n24) );
  NAND2_X1 U7 ( .A1(n29), .A2(n22), .ZN(n27) );
  INV_X1 U8 ( .A(n28), .ZN(n25) );
  OAI21_X1 U9 ( .B1(n20), .B2(n21), .A(n22), .ZN(n13) );
  OAI21_X1 U10 ( .B1(n20), .B2(n23), .A(n22), .ZN(n16) );
  AOI21_X1 U11 ( .B1(n16), .B2(n12), .A(n14), .ZN(n15) );
  AOI21_X1 U12 ( .B1(n12), .B2(n13), .A(n14), .ZN(n10) );
  AOI21_X1 U13 ( .B1(n23), .B2(n8), .A(n21), .ZN(n26) );
  OAI21_X1 U14 ( .B1(n8), .B2(n21), .A(n23), .ZN(n28) );
  INV_X1 U15 ( .A(n17), .ZN(n14) );
  INV_X1 U16 ( .A(n20), .ZN(n29) );
  XNOR2_X1 U17 ( .A(n15), .B(n11), .ZN(n7) );
  XNOR2_X1 U18 ( .A(n10), .B(n11), .ZN(n9) );
  XNOR2_X1 U19 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  NOR2_X1 U20 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  NAND2_X1 U21 ( .A1(B[0]), .A2(A[0]), .ZN(n23) );
  OR2_X1 U22 ( .A1(A[2]), .A2(B[2]), .ZN(n12) );
  NAND2_X1 U23 ( .A1(B[2]), .A2(A[2]), .ZN(n17) );
  OAI22_X1 U24 ( .A1(Ci), .A2(n7), .B1(n8), .B2(n9), .ZN(S[3]) );
  OAI21_X1 U25 ( .B1(Ci), .B2(n16), .A(n13), .ZN(n19) );
  INV_X1 U26 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n22) );
  NOR2_X1 U28 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
endmodule


module carry_sel_bk_NB4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  wire   n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32;

  XOR2_X1 U28 ( .A(n17), .B(n18), .Z(S[2]) );
  XOR2_X1 U29 ( .A(n32), .B(n29), .Z(S[0]) );
  NAND2_X1 U2 ( .A1(n30), .A2(n23), .ZN(n29) );
  INV_X1 U3 ( .A(n22), .ZN(n30) );
  OAI22_X1 U4 ( .A1(n31), .A2(n20), .B1(n21), .B2(n23), .ZN(n16) );
  OAI22_X1 U5 ( .A1(n31), .A2(n20), .B1(n21), .B2(n22), .ZN(n12) );
  OAI21_X1 U6 ( .B1(n12), .B2(n13), .A(n14), .ZN(n11) );
  OAI21_X1 U7 ( .B1(n32), .B2(n22), .A(n23), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n13), .B2(n16), .A(n14), .ZN(n15) );
  OAI22_X1 U9 ( .A1(n24), .A2(n25), .B1(n26), .B2(n27), .ZN(S[1]) );
  INV_X1 U10 ( .A(n28), .ZN(n26) );
  AOI21_X1 U11 ( .B1(n23), .B2(n32), .A(n22), .ZN(n24) );
  INV_X1 U12 ( .A(n27), .ZN(n25) );
  OAI21_X1 U13 ( .B1(Ci), .B2(n16), .A(n12), .ZN(n17) );
  OAI22_X1 U14 ( .A1(Ci), .A2(n7), .B1(n8), .B2(n32), .ZN(S[3]) );
  XNOR2_X1 U15 ( .A(n15), .B(n10), .ZN(n7) );
  XNOR2_X1 U16 ( .A(n10), .B(n11), .ZN(n8) );
  INV_X1 U17 ( .A(A[1]), .ZN(n31) );
  XNOR2_X1 U18 ( .A(n31), .B(B[1]), .ZN(n27) );
  INV_X1 U19 ( .A(B[1]), .ZN(n20) );
  NOR2_X1 U20 ( .A1(B[1]), .A2(A[1]), .ZN(n21) );
  XNOR2_X1 U21 ( .A(B[3]), .B(A[3]), .ZN(n10) );
  XNOR2_X1 U22 ( .A(A[2]), .B(B[2]), .ZN(n18) );
  AND2_X1 U23 ( .A1(B[2]), .A2(A[2]), .ZN(n13) );
  OR2_X1 U24 ( .A1(A[2]), .A2(B[2]), .ZN(n14) );
  NAND2_X1 U25 ( .A1(B[0]), .A2(A[0]), .ZN(n23) );
  NOR2_X1 U26 ( .A1(B[0]), .A2(A[0]), .ZN(n22) );
  INV_X1 U27 ( .A(Ci), .ZN(n32) );
endmodule


module G_76 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
endmodule


module G_77 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
endmodule


module blockPG_219 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module G_79 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
endmodule


module blockPG_230 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module blockPG_237 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
endmodule


module blockPG_241 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
endmodule


module G_0 ( Gik, Gk_1j, Pik, Gij );
  input Gik, Gk_1j, Pik;
  output Gij;
  wire   n2;

  AOI21_X1 U1 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(Gij) );
endmodule


module blockPG_0 ( Gik, Gk_1j, Pik, Pk_1j, Pij, Gij );
  input Gik, Gk_1j, Pik, Pk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
endmodule


module pg_net_260 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_263 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_285 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_287 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_0 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module p4addgen_NB32_CW4_1 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_1 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_1 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_2 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_2 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_2 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_3 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_3 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_3 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_4 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_4 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_4 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_5 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_5 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_5 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_6 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_6 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_6 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_7 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_7 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_7 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module p4addgen_NB32_CW4_8 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_8 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_8 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module MUX_SHIFT_NB16_N_sh14 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   \B[30] , AS, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n46,
         \B[6] , \B[1] , \B[12] , n97;
  assign B[31] = \B[30] ;
  assign B[30] = \B[30] ;
  assign B[5] = AS;
  assign B[10] = \B[6] ;
  assign B[13] = \B[6] ;
  assign B[2] = \B[6] ;
  assign B[6] = \B[6] ;
  assign B[4] = \B[1] ;
  assign B[8] = \B[1] ;
  assign B[9] = \B[1] ;
  assign B[1] = \B[1] ;
  assign B[3] = \B[12] ;
  assign B[11] = \B[12] ;
  assign B[7] = \B[12] ;
  assign B[0] = \B[12] ;
  assign B[12] = \B[12] ;

  XOR2_X1 U30 ( .A(sel[1]), .B(A[14]), .Z(n13) );
  XOR2_X1 U31 ( .A(A[15]), .B(n9), .Z(n7) );
  XOR2_X1 U32 ( .A(sel[1]), .B(A[13]), .Z(n15) );
  XOR2_X1 U33 ( .A(A[14]), .B(n9), .Z(n14) );
  XOR2_X1 U34 ( .A(sel[1]), .B(A[12]), .Z(n17) );
  XOR2_X1 U35 ( .A(A[13]), .B(n9), .Z(n16) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[11]), .Z(n19) );
  XOR2_X1 U37 ( .A(A[12]), .B(n9), .Z(n18) );
  XOR2_X1 U38 ( .A(sel[1]), .B(A[10]), .Z(n21) );
  XOR2_X1 U39 ( .A(A[11]), .B(n9), .Z(n20) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[9]), .Z(n23) );
  XOR2_X1 U41 ( .A(A[10]), .B(n9), .Z(n22) );
  XOR2_X1 U42 ( .A(sel[1]), .B(A[8]), .Z(n25) );
  XOR2_X1 U43 ( .A(A[9]), .B(n9), .Z(n24) );
  XOR2_X1 U44 ( .A(sel[1]), .B(A[7]), .Z(n27) );
  XOR2_X1 U45 ( .A(A[8]), .B(n9), .Z(n26) );
  XOR2_X1 U46 ( .A(sel[1]), .B(A[6]), .Z(n29) );
  XOR2_X1 U47 ( .A(A[7]), .B(n9), .Z(n28) );
  XOR2_X1 U48 ( .A(sel[1]), .B(A[5]), .Z(n31) );
  XOR2_X1 U49 ( .A(A[6]), .B(n9), .Z(n30) );
  XOR2_X1 U50 ( .A(sel[1]), .B(A[4]), .Z(n33) );
  XOR2_X1 U51 ( .A(A[5]), .B(n9), .Z(n32) );
  XOR2_X1 U52 ( .A(sel[1]), .B(A[3]), .Z(n35) );
  XOR2_X1 U53 ( .A(A[4]), .B(n9), .Z(n34) );
  XOR2_X1 U54 ( .A(sel[1]), .B(A[2]), .Z(n37) );
  XOR2_X1 U55 ( .A(A[3]), .B(n9), .Z(n36) );
  XOR2_X1 U56 ( .A(sel[1]), .B(A[1]), .Z(n39) );
  XOR2_X1 U57 ( .A(A[2]), .B(n9), .Z(n38) );
  XOR2_X1 U58 ( .A(sel[1]), .B(A[0]), .Z(n41) );
  XOR2_X1 U59 ( .A(n9), .B(n43), .Z(n42) );
  XOR2_X1 U60 ( .A(A[1]), .B(n9), .Z(n40) );
  XOR2_X1 U61 ( .A(sel[0]), .B(sel[1]), .Z(n10) );
  OAI21_X1 U3 ( .B1(n6), .B2(n7), .A(n8), .ZN(\B[30] ) );
  INV_X1 U4 ( .A(n10), .ZN(n11) );
  NAND2_X1 U5 ( .A1(n11), .A2(n42), .ZN(n12) );
  OAI22_X1 U6 ( .A1(n11), .A2(n26), .B1(n12), .B2(n27), .ZN(B[22]) );
  OAI22_X1 U7 ( .A1(n11), .A2(n34), .B1(n12), .B2(n35), .ZN(B[18]) );
  OAI22_X1 U8 ( .A1(n11), .A2(n18), .B1(n12), .B2(n19), .ZN(B[26]) );
  OAI22_X1 U9 ( .A1(n44), .A2(n97), .B1(sel[2]), .B2(n46), .ZN(B[14]) );
  INV_X1 U10 ( .A(n46), .ZN(n44) );
  OAI22_X1 U11 ( .A1(n11), .A2(n28), .B1(n12), .B2(n29), .ZN(B[21]) );
  OAI22_X1 U12 ( .A1(n11), .A2(n36), .B1(n12), .B2(n37), .ZN(B[17]) );
  OAI22_X1 U13 ( .A1(n11), .A2(n20), .B1(n12), .B2(n21), .ZN(B[25]) );
  OAI22_X1 U14 ( .A1(n11), .A2(n7), .B1(n12), .B2(n13), .ZN(B[29]) );
  OAI22_X1 U15 ( .A1(n11), .A2(n30), .B1(n12), .B2(n31), .ZN(B[20]) );
  OAI22_X1 U16 ( .A1(n11), .A2(n38), .B1(n12), .B2(n39), .ZN(B[16]) );
  OAI22_X1 U17 ( .A1(n11), .A2(n22), .B1(n12), .B2(n23), .ZN(B[24]) );
  OAI22_X1 U18 ( .A1(n11), .A2(n14), .B1(n12), .B2(n15), .ZN(B[28]) );
  OAI22_X1 U19 ( .A1(n11), .A2(n40), .B1(n12), .B2(n41), .ZN(B[15]) );
  OAI22_X1 U20 ( .A1(n11), .A2(n16), .B1(n12), .B2(n17), .ZN(B[27]) );
  OAI22_X1 U21 ( .A1(n11), .A2(n24), .B1(n12), .B2(n25), .ZN(B[23]) );
  OAI22_X1 U22 ( .A1(n11), .A2(n32), .B1(n12), .B2(n33), .ZN(B[19]) );
  INV_X1 U23 ( .A(sel[2]), .ZN(n9) );
  AOI21_X1 U24 ( .B1(sel[1]), .B2(A[15]), .A(n10), .ZN(n6) );
  AOI21_X1 U25 ( .B1(sel[1]), .B2(sel[0]), .A(n9), .ZN(AS) );
  INV_X1 U26 ( .A(sel[1]), .ZN(n43) );
  OR3_X1 U27 ( .A1(A[15]), .A2(sel[1]), .A3(n9), .ZN(n8) );
  NAND2_X1 U28 ( .A1(A[0]), .A2(n10), .ZN(n46) );
  INV_X1 U29 ( .A(n97), .ZN(\B[6] ) );
  INV_X1 U62 ( .A(n97), .ZN(\B[1] ) );
  INV_X1 U63 ( .A(n97), .ZN(\B[12] ) );
  INV_X1 U64 ( .A(AS), .ZN(n97) );
endmodule


module MUX_SHIFT_NB16_N_sh12 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   \B[7] , n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n46,
         \B[2] , \B[6] , \B[9] , n67;
  assign B[31] = B[28];
  assign B[30] = B[28];
  assign B[29] = B[28];
  assign B[11] = \B[7] ;
  assign B[3] = \B[7] ;
  assign B[7] = \B[7] ;
  assign B[5] = \B[2] ;
  assign B[10] = \B[2] ;
  assign B[2] = \B[2] ;
  assign B[1] = \B[6] ;
  assign AS = \B[6] ;
  assign B[6] = \B[6] ;
  assign B[0] = \B[9] ;
  assign B[4] = \B[9] ;
  assign B[8] = \B[9] ;
  assign B[9] = \B[9] ;

  OAI21_X2 U3 ( .B1(n6), .B2(n7), .A(n8), .ZN(B[28]) );
  XOR2_X1 U30 ( .A(sel[1]), .B(A[14]), .Z(n13) );
  XOR2_X1 U31 ( .A(A[15]), .B(n9), .Z(n7) );
  XOR2_X1 U32 ( .A(sel[1]), .B(A[13]), .Z(n15) );
  XOR2_X1 U33 ( .A(A[14]), .B(n9), .Z(n14) );
  XOR2_X1 U34 ( .A(sel[1]), .B(A[12]), .Z(n17) );
  XOR2_X1 U35 ( .A(A[13]), .B(n9), .Z(n16) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[11]), .Z(n19) );
  XOR2_X1 U37 ( .A(A[12]), .B(n9), .Z(n18) );
  XOR2_X1 U38 ( .A(sel[1]), .B(A[10]), .Z(n21) );
  XOR2_X1 U39 ( .A(A[11]), .B(n9), .Z(n20) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[9]), .Z(n23) );
  XOR2_X1 U41 ( .A(A[10]), .B(n9), .Z(n22) );
  XOR2_X1 U42 ( .A(sel[1]), .B(A[8]), .Z(n25) );
  XOR2_X1 U43 ( .A(A[9]), .B(n9), .Z(n24) );
  XOR2_X1 U44 ( .A(sel[1]), .B(A[7]), .Z(n27) );
  XOR2_X1 U45 ( .A(A[8]), .B(n9), .Z(n26) );
  XOR2_X1 U46 ( .A(sel[1]), .B(A[6]), .Z(n29) );
  XOR2_X1 U47 ( .A(A[7]), .B(n9), .Z(n28) );
  XOR2_X1 U48 ( .A(sel[1]), .B(A[5]), .Z(n31) );
  XOR2_X1 U49 ( .A(A[6]), .B(n9), .Z(n30) );
  XOR2_X1 U50 ( .A(sel[1]), .B(A[4]), .Z(n33) );
  XOR2_X1 U51 ( .A(A[5]), .B(n9), .Z(n32) );
  XOR2_X1 U52 ( .A(sel[1]), .B(A[3]), .Z(n35) );
  XOR2_X1 U53 ( .A(A[4]), .B(n9), .Z(n34) );
  XOR2_X1 U54 ( .A(sel[1]), .B(A[2]), .Z(n37) );
  XOR2_X1 U55 ( .A(A[3]), .B(n9), .Z(n36) );
  XOR2_X1 U56 ( .A(sel[1]), .B(A[1]), .Z(n39) );
  XOR2_X1 U57 ( .A(A[2]), .B(n9), .Z(n38) );
  XOR2_X1 U58 ( .A(sel[1]), .B(A[0]), .Z(n41) );
  XOR2_X1 U59 ( .A(n9), .B(n43), .Z(n42) );
  XOR2_X1 U60 ( .A(A[1]), .B(n9), .Z(n40) );
  XOR2_X1 U61 ( .A(sel[0]), .B(sel[1]), .Z(n10) );
  INV_X1 U4 ( .A(n10), .ZN(n11) );
  OR3_X1 U5 ( .A1(A[15]), .A2(sel[1]), .A3(n9), .ZN(n8) );
  AOI21_X1 U6 ( .B1(sel[1]), .B2(A[15]), .A(n10), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n11), .A2(n42), .ZN(n12) );
  INV_X1 U8 ( .A(sel[1]), .ZN(n43) );
  OAI22_X1 U9 ( .A1(n11), .A2(n38), .B1(n12), .B2(n39), .ZN(B[14]) );
  OAI22_X1 U10 ( .A1(n11), .A2(n14), .B1(n12), .B2(n15), .ZN(B[26]) );
  OAI22_X1 U11 ( .A1(n11), .A2(n30), .B1(n12), .B2(n31), .ZN(B[18]) );
  OAI22_X1 U12 ( .A1(n11), .A2(n22), .B1(n12), .B2(n23), .ZN(B[22]) );
  INV_X1 U13 ( .A(sel[2]), .ZN(n9) );
  OAI22_X1 U14 ( .A1(n11), .A2(n40), .B1(n12), .B2(n41), .ZN(B[13]) );
  OAI22_X1 U15 ( .A1(n11), .A2(n16), .B1(n12), .B2(n17), .ZN(B[25]) );
  OAI22_X1 U16 ( .A1(n11), .A2(n32), .B1(n12), .B2(n33), .ZN(B[17]) );
  OAI22_X1 U17 ( .A1(n11), .A2(n24), .B1(n12), .B2(n25), .ZN(B[21]) );
  OAI22_X1 U18 ( .A1(n11), .A2(n18), .B1(n12), .B2(n19), .ZN(B[24]) );
  OAI22_X1 U19 ( .A1(n11), .A2(n34), .B1(n12), .B2(n35), .ZN(B[16]) );
  OAI22_X1 U20 ( .A1(n11), .A2(n26), .B1(n12), .B2(n27), .ZN(B[20]) );
  OAI22_X1 U21 ( .A1(n44), .A2(n67), .B1(sel[2]), .B2(n46), .ZN(B[12]) );
  INV_X1 U22 ( .A(n46), .ZN(n44) );
  OAI22_X1 U23 ( .A1(n11), .A2(n7), .B1(n12), .B2(n13), .ZN(B[27]) );
  OAI22_X1 U24 ( .A1(n11), .A2(n36), .B1(n12), .B2(n37), .ZN(B[15]) );
  OAI22_X1 U25 ( .A1(n11), .A2(n28), .B1(n12), .B2(n29), .ZN(B[19]) );
  OAI22_X1 U26 ( .A1(n11), .A2(n20), .B1(n12), .B2(n21), .ZN(B[23]) );
  AOI21_X1 U27 ( .B1(sel[1]), .B2(sel[0]), .A(n9), .ZN(\B[7] ) );
  NAND2_X1 U28 ( .A1(A[0]), .A2(n10), .ZN(n46) );
  INV_X1 U29 ( .A(n67), .ZN(\B[2] ) );
  INV_X1 U62 ( .A(n67), .ZN(\B[6] ) );
  INV_X1 U63 ( .A(n67), .ZN(\B[9] ) );
  INV_X1 U64 ( .A(\B[7] ), .ZN(n67) );
endmodule


module MUX_SHIFT_NB16_N_sh10 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   n69, \B[5]_snps_wire , n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, \B[2] , AS, \B[4] ;
  assign B[31] = B[26];
  assign B[27] = B[26];
  assign B[28] = B[26];
  assign B[29] = B[26];
  assign B[30] = B[26];
  assign B[1] = \B[2] ;
  assign B[6] = \B[2] ;
  assign B[2] = \B[2] ;
  assign B[7] = AS;
  assign B[9] = AS;
  assign B[5] = AS;
  assign B[3] = \B[4] ;
  assign B[0] = \B[4] ;
  assign B[8] = \B[4] ;
  assign B[4] = \B[4] ;

  XOR2_X1 U30 ( .A(sel[1]), .B(A[14]), .Z(n13) );
  XOR2_X1 U31 ( .A(A[15]), .B(n9), .Z(n7) );
  XOR2_X1 U32 ( .A(sel[1]), .B(A[13]), .Z(n15) );
  XOR2_X1 U33 ( .A(A[14]), .B(n9), .Z(n14) );
  XOR2_X1 U34 ( .A(sel[1]), .B(A[12]), .Z(n17) );
  XOR2_X1 U35 ( .A(A[13]), .B(n9), .Z(n16) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[11]), .Z(n19) );
  XOR2_X1 U37 ( .A(A[12]), .B(n9), .Z(n18) );
  XOR2_X1 U38 ( .A(sel[1]), .B(A[10]), .Z(n21) );
  XOR2_X1 U39 ( .A(A[11]), .B(n9), .Z(n20) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[9]), .Z(n23) );
  XOR2_X1 U41 ( .A(A[10]), .B(n9), .Z(n22) );
  XOR2_X1 U42 ( .A(sel[1]), .B(A[8]), .Z(n25) );
  XOR2_X1 U43 ( .A(A[9]), .B(n9), .Z(n24) );
  XOR2_X1 U44 ( .A(sel[1]), .B(A[7]), .Z(n27) );
  XOR2_X1 U45 ( .A(A[8]), .B(n9), .Z(n26) );
  XOR2_X1 U46 ( .A(sel[1]), .B(A[6]), .Z(n29) );
  XOR2_X1 U47 ( .A(A[7]), .B(n9), .Z(n28) );
  XOR2_X1 U48 ( .A(sel[1]), .B(A[5]), .Z(n31) );
  XOR2_X1 U49 ( .A(A[6]), .B(n9), .Z(n30) );
  XOR2_X1 U50 ( .A(sel[1]), .B(A[4]), .Z(n33) );
  XOR2_X1 U51 ( .A(A[5]), .B(n9), .Z(n32) );
  XOR2_X1 U52 ( .A(sel[1]), .B(A[3]), .Z(n35) );
  XOR2_X1 U53 ( .A(A[4]), .B(n9), .Z(n34) );
  XOR2_X1 U54 ( .A(sel[1]), .B(A[2]), .Z(n37) );
  XOR2_X1 U55 ( .A(A[3]), .B(n9), .Z(n36) );
  XOR2_X1 U56 ( .A(sel[1]), .B(A[1]), .Z(n39) );
  XOR2_X1 U57 ( .A(A[2]), .B(n9), .Z(n38) );
  XOR2_X1 U58 ( .A(sel[1]), .B(A[0]), .Z(n41) );
  XOR2_X1 U59 ( .A(n9), .B(n43), .Z(n42) );
  XOR2_X1 U60 ( .A(A[1]), .B(n9), .Z(n40) );
  XOR2_X1 U61 ( .A(sel[0]), .B(sel[1]), .Z(n10) );
  INV_X1 U3 ( .A(n10), .ZN(n11) );
  BUF_X2 U4 ( .A(n69), .Z(B[26]) );
  OAI21_X1 U5 ( .B1(n6), .B2(n7), .A(n8), .ZN(n69) );
  OR3_X1 U6 ( .A1(A[15]), .A2(sel[1]), .A3(n9), .ZN(n8) );
  AOI21_X1 U7 ( .B1(A[15]), .B2(sel[1]), .A(n10), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n11), .A2(n42), .ZN(n12) );
  INV_X1 U9 ( .A(sel[1]), .ZN(n43) );
  OAI22_X1 U10 ( .A1(n11), .A2(n34), .B1(n12), .B2(n35), .ZN(B[14]) );
  OAI22_X1 U11 ( .A1(n11), .A2(n26), .B1(n12), .B2(n27), .ZN(B[18]) );
  OAI22_X1 U12 ( .A1(n11), .A2(n18), .B1(n12), .B2(n19), .ZN(B[22]) );
  OAI22_X1 U13 ( .A1(n11), .A2(n36), .B1(n12), .B2(n37), .ZN(B[13]) );
  OAI22_X1 U14 ( .A1(n11), .A2(n7), .B1(n12), .B2(n13), .ZN(B[25]) );
  OAI22_X1 U15 ( .A1(n11), .A2(n28), .B1(n12), .B2(n29), .ZN(B[17]) );
  OAI22_X1 U16 ( .A1(n11), .A2(n20), .B1(n12), .B2(n21), .ZN(B[21]) );
  OAI22_X1 U17 ( .A1(n11), .A2(n14), .B1(n12), .B2(n15), .ZN(B[24]) );
  OAI22_X1 U18 ( .A1(n11), .A2(n38), .B1(n12), .B2(n39), .ZN(B[12]) );
  OAI22_X1 U19 ( .A1(n11), .A2(n30), .B1(n12), .B2(n31), .ZN(B[16]) );
  OAI22_X1 U20 ( .A1(n11), .A2(n22), .B1(n12), .B2(n23), .ZN(B[20]) );
  OAI22_X1 U21 ( .A1(n11), .A2(n40), .B1(n12), .B2(n41), .ZN(B[11]) );
  OAI22_X1 U22 ( .A1(n11), .A2(n32), .B1(n12), .B2(n33), .ZN(B[15]) );
  OAI22_X1 U23 ( .A1(n11), .A2(n24), .B1(n12), .B2(n25), .ZN(B[19]) );
  OAI22_X1 U24 ( .A1(n11), .A2(n16), .B1(n12), .B2(n17), .ZN(B[23]) );
  INV_X1 U25 ( .A(sel[2]), .ZN(n9) );
  INV_X1 U26 ( .A(n44), .ZN(B[10]) );
  AOI22_X1 U27 ( .A1(n45), .A2(\B[4] ), .B1(n9), .B2(n46), .ZN(n44) );
  INV_X1 U28 ( .A(n45), .ZN(n46) );
  AOI21_X1 U29 ( .B1(sel[0]), .B2(sel[1]), .A(n9), .ZN(\B[5]_snps_wire ) );
  NAND2_X1 U62 ( .A1(A[0]), .A2(n10), .ZN(n45) );
  CLKBUF_X1 U63 ( .A(\B[5]_snps_wire ), .Z(\B[2] ) );
  CLKBUF_X1 U64 ( .A(\B[5]_snps_wire ), .Z(AS) );
  CLKBUF_X1 U65 ( .A(\B[5]_snps_wire ), .Z(\B[4] ) );
endmodule


module MUX_SHIFT_NB16_N_sh8 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_24, \B[1]_snps_wire , n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, \B[6] , \B[26] ;
  assign B[7] = \B[6] ;
  assign B[3] = \B[6] ;
  assign B[4] = \B[6] ;
  assign B[0] = \B[6] ;
  assign B[5] = \B[6] ;
  assign B[1] = \B[6] ;
  assign AS = \B[6] ;
  assign B[2] = \B[6] ;
  assign B[6] = \B[6] ;
  assign B[31] = \B[26] ;
  assign B[27] = \B[26] ;
  assign B[24] = \B[26] ;
  assign B[28] = \B[26] ;
  assign B[29] = \B[26] ;
  assign B[25] = \B[26] ;
  assign B[30] = \B[26] ;
  assign B[26] = \B[26] ;

  XOR2_X2 U3 ( .A(sel[0]), .B(n10), .Z(n6) );
  BUF_X2 U4 ( .A(\B[1]_snps_wire ), .Z(\B[6] ) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n10) );
  INV_X1 U6 ( .A(n6), .ZN(n15) );
  NAND2_X1 U7 ( .A1(n6), .A2(n46), .ZN(n8) );
  BUF_X2 U8 ( .A(B_24), .Z(\B[26] ) );
  OAI21_X1 U9 ( .B1(n16), .B2(n17), .A(n18), .ZN(B_24) );
  OR3_X1 U10 ( .A1(A[15]), .A2(sel[1]), .A3(n13), .ZN(n18) );
  AOI21_X1 U11 ( .B1(A[15]), .B2(sel[1]), .A(n15), .ZN(n16) );
  OAI22_X1 U12 ( .A1(n6), .A2(n44), .B1(n8), .B2(n45), .ZN(B[10]) );
  XNOR2_X1 U13 ( .A(n10), .B(A[1]), .ZN(n45) );
  OAI22_X1 U14 ( .A1(n6), .A2(n36), .B1(n8), .B2(n37), .ZN(B[14]) );
  OAI22_X1 U15 ( .A1(n6), .A2(n28), .B1(n8), .B2(n29), .ZN(B[18]) );
  XNOR2_X1 U16 ( .A(n10), .B(A[9]), .ZN(n29) );
  OAI22_X1 U17 ( .A1(n6), .A2(n20), .B1(n8), .B2(n21), .ZN(B[22]) );
  OAI22_X1 U18 ( .A1(n6), .A2(n7), .B1(n8), .B2(n9), .ZN(B[9]) );
  OAI22_X1 U19 ( .A1(n6), .A2(n38), .B1(n8), .B2(n39), .ZN(B[13]) );
  XNOR2_X1 U20 ( .A(n10), .B(A[4]), .ZN(n39) );
  OAI22_X1 U21 ( .A1(n6), .A2(n30), .B1(n8), .B2(n31), .ZN(B[17]) );
  XNOR2_X1 U22 ( .A(n10), .B(A[8]), .ZN(n31) );
  OAI22_X1 U23 ( .A1(n6), .A2(n22), .B1(n8), .B2(n23), .ZN(B[21]) );
  XNOR2_X1 U24 ( .A(n10), .B(A[12]), .ZN(n23) );
  OAI22_X1 U25 ( .A1(n6), .A2(n40), .B1(n8), .B2(n41), .ZN(B[12]) );
  XNOR2_X1 U26 ( .A(n10), .B(A[3]), .ZN(n41) );
  OAI22_X1 U27 ( .A1(n6), .A2(n32), .B1(n8), .B2(n33), .ZN(B[16]) );
  XNOR2_X1 U28 ( .A(n10), .B(A[7]), .ZN(n33) );
  OAI22_X1 U29 ( .A1(n6), .A2(n24), .B1(n8), .B2(n25), .ZN(B[20]) );
  XNOR2_X1 U30 ( .A(n10), .B(A[11]), .ZN(n25) );
  OAI22_X1 U31 ( .A1(n6), .A2(n42), .B1(n8), .B2(n43), .ZN(B[11]) );
  OAI22_X1 U32 ( .A1(n6), .A2(n34), .B1(n8), .B2(n35), .ZN(B[15]) );
  XNOR2_X1 U33 ( .A(n10), .B(A[6]), .ZN(n35) );
  OAI22_X1 U34 ( .A1(n6), .A2(n26), .B1(n8), .B2(n27), .ZN(B[19]) );
  XNOR2_X1 U35 ( .A(n10), .B(A[10]), .ZN(n27) );
  OAI22_X1 U36 ( .A1(n6), .A2(n17), .B1(n8), .B2(n19), .ZN(B[23]) );
  XNOR2_X1 U37 ( .A(n10), .B(A[14]), .ZN(n19) );
  AOI21_X1 U38 ( .B1(sel[1]), .B2(sel[0]), .A(n13), .ZN(\B[1]_snps_wire ) );
  INV_X1 U39 ( .A(n11), .ZN(B[8]) );
  AOI22_X1 U40 ( .A1(n12), .A2(\B[6] ), .B1(n13), .B2(n14), .ZN(n11) );
  INV_X1 U41 ( .A(n12), .ZN(n14) );
  XNOR2_X1 U42 ( .A(n10), .B(A[13]), .ZN(n21) );
  XNOR2_X1 U43 ( .A(n10), .B(A[2]), .ZN(n43) );
  XNOR2_X1 U44 ( .A(n10), .B(A[5]), .ZN(n37) );
  INV_X1 U45 ( .A(sel[2]), .ZN(n13) );
  XNOR2_X1 U46 ( .A(sel[2]), .B(n10), .ZN(n46) );
  XNOR2_X1 U47 ( .A(A[3]), .B(sel[2]), .ZN(n42) );
  XNOR2_X1 U48 ( .A(A[2]), .B(sel[2]), .ZN(n44) );
  XNOR2_X1 U49 ( .A(A[5]), .B(sel[2]), .ZN(n38) );
  XNOR2_X1 U50 ( .A(A[6]), .B(sel[2]), .ZN(n36) );
  XNOR2_X1 U51 ( .A(A[4]), .B(sel[2]), .ZN(n40) );
  XNOR2_X1 U52 ( .A(A[15]), .B(sel[2]), .ZN(n17) );
  XNOR2_X1 U53 ( .A(A[14]), .B(sel[2]), .ZN(n20) );
  XNOR2_X1 U54 ( .A(A[10]), .B(sel[2]), .ZN(n28) );
  XNOR2_X1 U55 ( .A(A[13]), .B(sel[2]), .ZN(n22) );
  XNOR2_X1 U56 ( .A(A[1]), .B(sel[2]), .ZN(n7) );
  XNOR2_X1 U57 ( .A(A[12]), .B(sel[2]), .ZN(n24) );
  XNOR2_X1 U58 ( .A(A[11]), .B(sel[2]), .ZN(n26) );
  XNOR2_X1 U59 ( .A(A[9]), .B(sel[2]), .ZN(n30) );
  XNOR2_X1 U60 ( .A(A[8]), .B(sel[2]), .ZN(n32) );
  XNOR2_X1 U61 ( .A(A[7]), .B(sel[2]), .ZN(n34) );
  NAND2_X1 U62 ( .A1(A[0]), .A2(n15), .ZN(n12) );
  XNOR2_X1 U63 ( .A(n10), .B(A[0]), .ZN(n9) );
endmodule


module MUX_SHIFT_NB16_N_sh6 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_24, AS, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n19, n20,
         n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         \B[1] , n65, \B[22] , \B[25] , n68, n69;
  assign B[5] = AS;
  assign B[2] = \B[1] ;
  assign B[3] = \B[1] ;
  assign B[0] = \B[1] ;
  assign B[4] = \B[1] ;
  assign B[1] = \B[1] ;
  assign B[27] = \B[22] ;
  assign B[29] = \B[22] ;
  assign B[26] = \B[22] ;
  assign B[30] = \B[22] ;
  assign B[22] = \B[22] ;
  assign B[31] = \B[25] ;
  assign B[23] = \B[25] ;
  assign B[28] = \B[25] ;
  assign B[24] = \B[25] ;
  assign B[25] = \B[25] ;

  XOR2_X1 U34 ( .A(sel[1]), .B(A[2]), .Z(n10) );
  XOR2_X1 U35 ( .A(A[3]), .B(n11), .Z(n8) );
  XOR2_X1 U36 ( .A(sel[1]), .B(A[1]), .Z(n13) );
  XOR2_X1 U37 ( .A(A[2]), .B(n11), .Z(n12) );
  XOR2_X1 U38 ( .A(A[1]), .B(n11), .Z(n14) );
  NAND3_X1 U39 ( .A1(sel[1]), .A2(n68), .A3(sel[0]), .ZN(n20) );
  XOR2_X1 U40 ( .A(sel[1]), .B(A[14]), .Z(n26) );
  XOR2_X1 U41 ( .A(sel[1]), .B(A[13]), .Z(n28) );
  XOR2_X1 U42 ( .A(A[14]), .B(n11), .Z(n27) );
  XOR2_X1 U43 ( .A(sel[1]), .B(A[12]), .Z(n30) );
  XOR2_X1 U44 ( .A(A[13]), .B(n11), .Z(n29) );
  XOR2_X1 U45 ( .A(sel[1]), .B(A[11]), .Z(n32) );
  XOR2_X1 U46 ( .A(A[12]), .B(n11), .Z(n31) );
  XOR2_X1 U47 ( .A(sel[1]), .B(A[10]), .Z(n34) );
  XOR2_X1 U48 ( .A(A[11]), .B(n11), .Z(n33) );
  XOR2_X1 U49 ( .A(sel[1]), .B(A[9]), .Z(n36) );
  XOR2_X1 U50 ( .A(A[10]), .B(n11), .Z(n35) );
  XOR2_X1 U51 ( .A(sel[1]), .B(A[8]), .Z(n38) );
  XOR2_X1 U52 ( .A(A[9]), .B(n11), .Z(n37) );
  XOR2_X1 U53 ( .A(sel[1]), .B(A[7]), .Z(n40) );
  XOR2_X1 U54 ( .A(A[8]), .B(n11), .Z(n39) );
  XOR2_X1 U55 ( .A(sel[1]), .B(A[6]), .Z(n42) );
  XOR2_X1 U56 ( .A(A[7]), .B(n11), .Z(n41) );
  XOR2_X1 U57 ( .A(sel[1]), .B(A[5]), .Z(n44) );
  XOR2_X1 U58 ( .A(A[6]), .B(n11), .Z(n43) );
  XOR2_X1 U59 ( .A(sel[1]), .B(A[4]), .Z(n46) );
  XOR2_X1 U60 ( .A(A[5]), .B(n11), .Z(n45) );
  XOR2_X1 U61 ( .A(sel[1]), .B(A[3]), .Z(n48) );
  XOR2_X1 U62 ( .A(sel[2]), .B(sel[1]), .Z(n49) );
  XOR2_X1 U63 ( .A(A[4]), .B(n11), .Z(n47) );
  XNOR2_X2 U3 ( .A(sel[0]), .B(sel[1]), .ZN(n7) );
  BUF_X1 U4 ( .A(B_24), .Z(\B[25] ) );
  NAND2_X1 U5 ( .A1(n7), .A2(n49), .ZN(n9) );
  OAI22_X1 U6 ( .A1(n7), .A2(n47), .B1(n9), .B2(n48), .ZN(B[10]) );
  OAI22_X1 U7 ( .A1(n7), .A2(n39), .B1(n9), .B2(n40), .ZN(B[14]) );
  OAI22_X1 U8 ( .A1(n7), .A2(n31), .B1(n9), .B2(n32), .ZN(B[18]) );
  OAI22_X1 U9 ( .A1(n7), .A2(n8), .B1(n9), .B2(n10), .ZN(B[9]) );
  OAI22_X1 U10 ( .A1(n7), .A2(n41), .B1(n9), .B2(n42), .ZN(B[13]) );
  OAI22_X1 U11 ( .A1(n7), .A2(n33), .B1(n9), .B2(n34), .ZN(B[17]) );
  OAI22_X1 U12 ( .A1(n7), .A2(n25), .B1(n9), .B2(n26), .ZN(B[21]) );
  INV_X1 U13 ( .A(n23), .ZN(n25) );
  OAI22_X1 U14 ( .A1(n7), .A2(n12), .B1(n9), .B2(n13), .ZN(B[8]) );
  OAI22_X1 U15 ( .A1(n7), .A2(n43), .B1(n9), .B2(n44), .ZN(B[12]) );
  OAI22_X1 U16 ( .A1(n7), .A2(n35), .B1(n9), .B2(n36), .ZN(B[16]) );
  OAI22_X1 U17 ( .A1(n7), .A2(n27), .B1(n9), .B2(n28), .ZN(B[20]) );
  OAI22_X1 U18 ( .A1(n17), .A2(n65), .B1(sel[2]), .B2(n19), .ZN(B[6]) );
  INV_X1 U19 ( .A(n17), .ZN(n19) );
  NOR2_X1 U20 ( .A1(n69), .A2(n7), .ZN(n17) );
  OAI22_X1 U21 ( .A1(n7), .A2(n45), .B1(n9), .B2(n46), .ZN(B[11]) );
  OAI22_X1 U22 ( .A1(n7), .A2(n37), .B1(n9), .B2(n38), .ZN(B[15]) );
  OAI22_X1 U23 ( .A1(n7), .A2(n14), .B1(n9), .B2(n15), .ZN(B[7]) );
  OAI22_X1 U24 ( .A1(n7), .A2(n29), .B1(n9), .B2(n30), .ZN(B[19]) );
  INV_X1 U25 ( .A(sel[2]), .ZN(n11) );
  XNOR2_X1 U26 ( .A(n68), .B(sel[2]), .ZN(n23) );
  AND2_X1 U27 ( .A1(n20), .A2(n21), .ZN(B_24) );
  OAI21_X1 U28 ( .B1(A[15]), .B2(n11), .A(n22), .ZN(n21) );
  OAI21_X1 U29 ( .B1(sel[1]), .B2(sel[0]), .A(n23), .ZN(n22) );
  AOI21_X1 U30 ( .B1(sel[1]), .B2(sel[0]), .A(n11), .ZN(AS) );
  XNOR2_X1 U31 ( .A(sel[1]), .B(n69), .ZN(n15) );
  INV_X1 U32 ( .A(n65), .ZN(\B[1] ) );
  INV_X1 U33 ( .A(AS), .ZN(n65) );
  CLKBUF_X2 U64 ( .A(B_24), .Z(\B[22] ) );
  INV_X1 U65 ( .A(A[15]), .ZN(n68) );
  INV_X1 U66 ( .A(A[0]), .ZN(n69) );
endmodule


module MUX_SHIFT_NB16_N_sh4 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   n70, \B[1]_snps_wire , n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, \B[2] , \B[22] , n68, n69;
  assign B[31] = B[21];
  assign B[23] = B[21];
  assign B[20] = B[21];
  assign B[24] = B[21];
  assign B[28] = B[21];
  assign B[29] = B[21];
  assign B[3] = \B[2] ;
  assign B[0] = \B[2] ;
  assign B[1] = \B[2] ;
  assign AS = \B[2] ;
  assign B[2] = \B[2] ;
  assign B[27] = \B[22] ;
  assign B[25] = \B[22] ;
  assign B[26] = \B[22] ;
  assign B[30] = \B[22] ;
  assign B[22] = \B[22] ;

  XOR2_X2 U3 ( .A(sel[0]), .B(n10), .Z(n6) );
  BUF_X1 U4 ( .A(\B[1]_snps_wire ), .Z(\B[2] ) );
  NAND2_X1 U5 ( .A1(n6), .A2(n46), .ZN(n8) );
  XNOR2_X1 U6 ( .A(n68), .B(n10), .ZN(n46) );
  INV_X1 U7 ( .A(n6), .ZN(n23) );
  XNOR2_X1 U8 ( .A(A[15]), .B(n68), .ZN(n25) );
  INV_X1 U9 ( .A(sel[1]), .ZN(n10) );
  OAI22_X1 U10 ( .A1(n6), .A2(n44), .B1(n8), .B2(n45), .ZN(B[10]) );
  XNOR2_X1 U11 ( .A(A[6]), .B(n68), .ZN(n44) );
  OAI22_X1 U12 ( .A1(n6), .A2(n36), .B1(n8), .B2(n37), .ZN(B[14]) );
  XNOR2_X1 U13 ( .A(A[10]), .B(n68), .ZN(n36) );
  XNOR2_X1 U14 ( .A(n10), .B(A[9]), .ZN(n37) );
  OAI22_X1 U15 ( .A1(n6), .A2(n28), .B1(n8), .B2(n29), .ZN(B[18]) );
  XNOR2_X1 U16 ( .A(A[14]), .B(n68), .ZN(n28) );
  OAI22_X1 U17 ( .A1(n6), .A2(n15), .B1(n8), .B2(n16), .ZN(B[6]) );
  XNOR2_X1 U18 ( .A(n10), .B(A[1]), .ZN(n16) );
  OAI22_X1 U19 ( .A1(n6), .A2(n7), .B1(n8), .B2(n9), .ZN(B[9]) );
  XNOR2_X1 U20 ( .A(n10), .B(A[4]), .ZN(n9) );
  OAI22_X1 U21 ( .A1(n6), .A2(n30), .B1(n8), .B2(n31), .ZN(B[17]) );
  XNOR2_X1 U22 ( .A(n10), .B(A[12]), .ZN(n31) );
  OAI22_X1 U23 ( .A1(n6), .A2(n17), .B1(n8), .B2(n18), .ZN(B[5]) );
  XNOR2_X1 U24 ( .A(A[1]), .B(n68), .ZN(n17) );
  OAI22_X1 U25 ( .A1(n6), .A2(n38), .B1(n8), .B2(n39), .ZN(B[13]) );
  XNOR2_X1 U26 ( .A(A[9]), .B(sel[2]), .ZN(n38) );
  XNOR2_X1 U27 ( .A(n10), .B(A[8]), .ZN(n39) );
  OAI22_X1 U28 ( .A1(n6), .A2(n11), .B1(n8), .B2(n12), .ZN(B[8]) );
  XNOR2_X1 U29 ( .A(n10), .B(A[3]), .ZN(n12) );
  XNOR2_X1 U30 ( .A(A[4]), .B(n68), .ZN(n11) );
  OAI22_X1 U31 ( .A1(n6), .A2(n32), .B1(n8), .B2(n33), .ZN(B[16]) );
  XNOR2_X1 U32 ( .A(n10), .B(A[11]), .ZN(n33) );
  XNOR2_X1 U33 ( .A(A[12]), .B(n68), .ZN(n32) );
  OAI22_X1 U34 ( .A1(n6), .A2(n40), .B1(n8), .B2(n41), .ZN(B[12]) );
  XNOR2_X1 U35 ( .A(A[8]), .B(sel[2]), .ZN(n40) );
  XNOR2_X1 U36 ( .A(n10), .B(A[7]), .ZN(n41) );
  OAI22_X1 U37 ( .A1(n6), .A2(n42), .B1(n8), .B2(n43), .ZN(B[11]) );
  XNOR2_X1 U38 ( .A(A[7]), .B(sel[2]), .ZN(n42) );
  XNOR2_X1 U39 ( .A(n10), .B(A[6]), .ZN(n43) );
  OAI22_X1 U40 ( .A1(n6), .A2(n34), .B1(n8), .B2(n35), .ZN(B[15]) );
  XNOR2_X1 U41 ( .A(A[11]), .B(n68), .ZN(n34) );
  XNOR2_X1 U42 ( .A(n10), .B(A[10]), .ZN(n35) );
  OAI22_X1 U43 ( .A1(n6), .A2(n25), .B1(n8), .B2(n27), .ZN(B[19]) );
  XNOR2_X1 U44 ( .A(n10), .B(A[14]), .ZN(n27) );
  OAI22_X1 U45 ( .A1(n6), .A2(n13), .B1(n8), .B2(n14), .ZN(B[7]) );
  XNOR2_X1 U46 ( .A(A[3]), .B(n68), .ZN(n13) );
  AOI21_X1 U47 ( .B1(sel[1]), .B2(sel[0]), .A(n69), .ZN(\B[1]_snps_wire ) );
  OAI21_X1 U48 ( .B1(n24), .B2(n25), .A(n26), .ZN(n70) );
  OR3_X1 U49 ( .A1(A[15]), .A2(sel[1]), .A3(n69), .ZN(n26) );
  AOI21_X1 U50 ( .B1(A[15]), .B2(sel[1]), .A(n23), .ZN(n24) );
  INV_X1 U51 ( .A(n19), .ZN(B[4]) );
  AOI22_X1 U52 ( .A1(n20), .A2(\B[2] ), .B1(n69), .B2(n22), .ZN(n19) );
  INV_X1 U53 ( .A(n20), .ZN(n22) );
  INV_X1 U54 ( .A(sel[2]), .ZN(n69) );
  XNOR2_X1 U55 ( .A(A[13]), .B(sel[2]), .ZN(n30) );
  XNOR2_X1 U56 ( .A(n10), .B(A[13]), .ZN(n29) );
  XNOR2_X1 U57 ( .A(A[2]), .B(n68), .ZN(n15) );
  XNOR2_X1 U58 ( .A(n10), .B(A[2]), .ZN(n14) );
  XNOR2_X1 U59 ( .A(A[5]), .B(sel[2]), .ZN(n7) );
  XNOR2_X1 U60 ( .A(n10), .B(A[5]), .ZN(n45) );
  NAND2_X1 U61 ( .A1(A[0]), .A2(n23), .ZN(n20) );
  XNOR2_X1 U62 ( .A(n10), .B(A[0]), .ZN(n18) );
  CLKBUF_X2 U63 ( .A(n70), .Z(\B[22] ) );
  CLKBUF_X2 U64 ( .A(n70), .Z(B[21]) );
  INV_X1 U65 ( .A(n69), .ZN(n68) );
endmodule


module MUX_SHIFT_NB16_N_sh2 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   \B[19]_snps_int_wire , \B[0] , n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, \B[30] , \B[24] , n66, n67;
  assign AS = \B[0] ;
  assign B[1] = \B[0] ;
  assign B[0] = \B[0] ;
  assign B[29] = \B[30] ;
  assign B[25] = \B[30] ;
  assign B[21] = \B[30] ;
  assign B[26] = \B[30] ;
  assign B[22] = \B[30] ;
  assign B[18] = \B[30] ;
  assign B[30] = \B[30] ;
  assign B[31] = \B[24] ;
  assign B[19] = \B[24] ;
  assign B[27] = \B[24] ;
  assign B[23] = \B[24] ;
  assign B[20] = \B[24] ;
  assign B[28] = \B[24] ;
  assign B[24] = \B[24] ;

  AOI21_X2 U59 ( .B1(sel[1]), .B2(sel[0]), .A(n67), .ZN(\B[0] ) );
  XOR2_X2 U3 ( .A(sel[0]), .B(n10), .Z(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(n46), .ZN(n8) );
  XNOR2_X1 U5 ( .A(n66), .B(n10), .ZN(n46) );
  BUF_X2 U6 ( .A(\B[19]_snps_int_wire ), .Z(\B[30] ) );
  BUF_X1 U7 ( .A(\B[19]_snps_int_wire ), .Z(\B[24] ) );
  INV_X1 U8 ( .A(n6), .ZN(n27) );
  XNOR2_X1 U9 ( .A(A[15]), .B(n66), .ZN(n29) );
  INV_X1 U10 ( .A(sel[1]), .ZN(n10) );
  OAI22_X1 U11 ( .A1(n6), .A2(n44), .B1(n8), .B2(n45), .ZN(B[10]) );
  XNOR2_X1 U12 ( .A(A[8]), .B(n66), .ZN(n44) );
  XNOR2_X1 U13 ( .A(n10), .B(A[7]), .ZN(n45) );
  OAI22_X1 U14 ( .A1(n6), .A2(n36), .B1(n8), .B2(n37), .ZN(B[14]) );
  XNOR2_X1 U15 ( .A(n10), .B(A[11]), .ZN(n37) );
  XNOR2_X1 U16 ( .A(A[12]), .B(sel[2]), .ZN(n36) );
  OAI22_X1 U17 ( .A1(n6), .A2(n15), .B1(n8), .B2(n16), .ZN(B[6]) );
  XNOR2_X1 U18 ( .A(n10), .B(A[3]), .ZN(n16) );
  XNOR2_X1 U19 ( .A(A[4]), .B(n66), .ZN(n15) );
  OAI22_X1 U20 ( .A1(n6), .A2(n7), .B1(n8), .B2(n9), .ZN(B[9]) );
  XNOR2_X1 U21 ( .A(A[7]), .B(n66), .ZN(n7) );
  XNOR2_X1 U22 ( .A(n10), .B(A[6]), .ZN(n9) );
  OAI22_X1 U23 ( .A1(n6), .A2(n17), .B1(n8), .B2(n18), .ZN(B[5]) );
  XNOR2_X1 U24 ( .A(A[3]), .B(n66), .ZN(n17) );
  OAI22_X1 U25 ( .A1(n6), .A2(n38), .B1(n8), .B2(n39), .ZN(B[13]) );
  XNOR2_X1 U26 ( .A(A[11]), .B(sel[2]), .ZN(n38) );
  XNOR2_X1 U27 ( .A(n10), .B(A[10]), .ZN(n39) );
  OAI22_X1 U28 ( .A1(n6), .A2(n29), .B1(n8), .B2(n31), .ZN(B[17]) );
  XNOR2_X1 U29 ( .A(n10), .B(A[14]), .ZN(n31) );
  OAI22_X1 U30 ( .A1(n6), .A2(n11), .B1(n8), .B2(n12), .ZN(B[8]) );
  XNOR2_X1 U31 ( .A(A[6]), .B(n66), .ZN(n11) );
  OAI22_X1 U32 ( .A1(n6), .A2(n19), .B1(n8), .B2(n20), .ZN(B[4]) );
  XNOR2_X1 U33 ( .A(n10), .B(A[1]), .ZN(n20) );
  OAI22_X1 U34 ( .A1(n6), .A2(n40), .B1(n8), .B2(n41), .ZN(B[12]) );
  XNOR2_X1 U35 ( .A(A[10]), .B(n66), .ZN(n40) );
  XNOR2_X1 U36 ( .A(n10), .B(A[9]), .ZN(n41) );
  OAI22_X1 U37 ( .A1(n6), .A2(n32), .B1(n8), .B2(n33), .ZN(B[16]) );
  XNOR2_X1 U38 ( .A(A[14]), .B(sel[2]), .ZN(n32) );
  OAI22_X1 U39 ( .A1(n6), .A2(n42), .B1(n8), .B2(n43), .ZN(B[11]) );
  XNOR2_X1 U40 ( .A(A[9]), .B(sel[2]), .ZN(n42) );
  XNOR2_X1 U41 ( .A(n10), .B(A[8]), .ZN(n43) );
  OAI22_X1 U42 ( .A1(n6), .A2(n34), .B1(n8), .B2(n35), .ZN(B[15]) );
  XNOR2_X1 U43 ( .A(n10), .B(A[12]), .ZN(n35) );
  OAI22_X1 U44 ( .A1(n6), .A2(n13), .B1(n8), .B2(n14), .ZN(B[7]) );
  XNOR2_X1 U45 ( .A(n10), .B(A[4]), .ZN(n14) );
  OAI22_X1 U46 ( .A1(n6), .A2(n21), .B1(n8), .B2(n22), .ZN(B[3]) );
  XNOR2_X1 U47 ( .A(A[1]), .B(n66), .ZN(n21) );
  INV_X1 U48 ( .A(n23), .ZN(B[2]) );
  AOI22_X1 U49 ( .A1(n24), .A2(\B[0] ), .B1(n67), .B2(n26), .ZN(n23) );
  INV_X1 U50 ( .A(n24), .ZN(n26) );
  OAI21_X1 U51 ( .B1(n28), .B2(n29), .A(n30), .ZN(\B[19]_snps_int_wire ) );
  OR3_X1 U52 ( .A1(A[15]), .A2(sel[1]), .A3(n67), .ZN(n30) );
  AOI21_X1 U53 ( .B1(A[15]), .B2(sel[1]), .A(n27), .ZN(n28) );
  INV_X1 U54 ( .A(sel[2]), .ZN(n67) );
  XNOR2_X1 U55 ( .A(A[13]), .B(sel[2]), .ZN(n34) );
  XNOR2_X1 U56 ( .A(n10), .B(A[13]), .ZN(n33) );
  XNOR2_X1 U57 ( .A(A[2]), .B(n66), .ZN(n19) );
  XNOR2_X1 U58 ( .A(n10), .B(A[2]), .ZN(n18) );
  XNOR2_X1 U60 ( .A(A[5]), .B(n66), .ZN(n13) );
  XNOR2_X1 U61 ( .A(n10), .B(A[5]), .ZN(n12) );
  NAND2_X1 U62 ( .A1(A[0]), .A2(n27), .ZN(n24) );
  XNOR2_X1 U63 ( .A(n10), .B(A[0]), .ZN(n22) );
  INV_X1 U64 ( .A(n67), .ZN(n66) );
endmodule


module MUX_SHIFT_NB16_N_sh0 ( A, sel, AS, B );
  input [15:0] A;
  input [2:0] sel;
  output [31:0] B;
  output AS;
  wire   B_17, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n45, n46,
         \B[30] , \B[29] , n67, n68, n69;
  assign B[21] = \B[30] ;
  assign B[25] = \B[30] ;
  assign B[17] = \B[30] ;
  assign B[22] = \B[30] ;
  assign B[18] = \B[30] ;
  assign B[26] = \B[30] ;
  assign B[30] = \B[30] ;
  assign B[31] = \B[29] ;
  assign B[27] = \B[29] ;
  assign B[19] = \B[29] ;
  assign B[23] = \B[29] ;
  assign B[28] = \B[29] ;
  assign B[24] = \B[29] ;
  assign B[16] = \B[29] ;
  assign B[20] = \B[29] ;
  assign B[29] = \B[29] ;

  XOR2_X1 U30 ( .A(n67), .B(A[8]), .Z(n9) );
  XOR2_X1 U31 ( .A(A[9]), .B(n10), .Z(n7) );
  XOR2_X1 U32 ( .A(n68), .B(A[7]), .Z(n12) );
  XOR2_X1 U33 ( .A(A[8]), .B(n10), .Z(n11) );
  XOR2_X1 U34 ( .A(n68), .B(A[6]), .Z(n14) );
  XOR2_X1 U35 ( .A(A[7]), .B(n10), .Z(n13) );
  XOR2_X1 U36 ( .A(n68), .B(A[5]), .Z(n16) );
  XOR2_X1 U37 ( .A(A[6]), .B(n10), .Z(n15) );
  XOR2_X1 U38 ( .A(n67), .B(A[4]), .Z(n18) );
  XOR2_X1 U39 ( .A(A[5]), .B(n10), .Z(n17) );
  XOR2_X1 U40 ( .A(n67), .B(A[3]), .Z(n20) );
  XOR2_X1 U41 ( .A(A[4]), .B(n10), .Z(n19) );
  XOR2_X1 U42 ( .A(n67), .B(A[2]), .Z(n22) );
  XOR2_X1 U43 ( .A(A[3]), .B(n10), .Z(n21) );
  XOR2_X1 U44 ( .A(n67), .B(A[1]), .Z(n24) );
  XOR2_X1 U45 ( .A(A[2]), .B(n10), .Z(n23) );
  XOR2_X1 U46 ( .A(n67), .B(A[0]), .Z(n26) );
  XOR2_X1 U47 ( .A(A[1]), .B(n10), .Z(n25) );
  XOR2_X1 U48 ( .A(n67), .B(A[14]), .Z(n31) );
  XOR2_X1 U49 ( .A(A[15]), .B(n10), .Z(n28) );
  XOR2_X1 U50 ( .A(n67), .B(A[13]), .Z(n33) );
  XOR2_X1 U51 ( .A(A[14]), .B(n10), .Z(n32) );
  XOR2_X1 U52 ( .A(n67), .B(A[12]), .Z(n35) );
  XOR2_X1 U53 ( .A(A[13]), .B(n10), .Z(n34) );
  XOR2_X1 U54 ( .A(n67), .B(A[11]), .Z(n37) );
  XOR2_X1 U55 ( .A(A[12]), .B(n10), .Z(n36) );
  XOR2_X1 U56 ( .A(n67), .B(A[10]), .Z(n39) );
  XOR2_X1 U57 ( .A(A[11]), .B(n10), .Z(n38) );
  XOR2_X1 U58 ( .A(n67), .B(A[9]), .Z(n41) );
  XOR2_X1 U59 ( .A(n10), .B(n69), .Z(n42) );
  XOR2_X1 U60 ( .A(A[10]), .B(n10), .Z(n40) );
  XOR2_X1 U61 ( .A(sel[0]), .B(n67), .Z(n30) );
  BUF_X2 U3 ( .A(B_17), .Z(\B[30] ) );
  NAND2_X1 U4 ( .A1(n6), .A2(n42), .ZN(n8) );
  BUF_X2 U5 ( .A(B_17), .Z(\B[29] ) );
  INV_X1 U6 ( .A(n69), .ZN(n67) );
  INV_X1 U7 ( .A(n30), .ZN(n6) );
  OAI22_X1 U8 ( .A1(n6), .A2(n40), .B1(n8), .B2(n41), .ZN(B[10]) );
  OAI22_X1 U9 ( .A1(n6), .A2(n15), .B1(n8), .B2(n16), .ZN(B[6]) );
  OAI22_X1 U10 ( .A1(n6), .A2(n32), .B1(n8), .B2(n33), .ZN(B[14]) );
  OAI22_X1 U11 ( .A1(n6), .A2(n23), .B1(n8), .B2(n24), .ZN(B[2]) );
  INV_X1 U12 ( .A(sel[2]), .ZN(n10) );
  OAI22_X1 U13 ( .A1(n6), .A2(n7), .B1(n8), .B2(n9), .ZN(B[9]) );
  OAI22_X1 U14 ( .A1(n6), .A2(n34), .B1(n8), .B2(n35), .ZN(B[13]) );
  OAI22_X1 U15 ( .A1(n6), .A2(n25), .B1(n8), .B2(n26), .ZN(B[1]) );
  OAI22_X1 U16 ( .A1(n6), .A2(n17), .B1(n8), .B2(n18), .ZN(B[5]) );
  OAI22_X1 U17 ( .A1(n6), .A2(n11), .B1(n8), .B2(n12), .ZN(B[8]) );
  OAI22_X1 U18 ( .A1(n6), .A2(n36), .B1(n8), .B2(n37), .ZN(B[12]) );
  OAI22_X1 U19 ( .A1(n6), .A2(n19), .B1(n8), .B2(n20), .ZN(B[4]) );
  OAI22_X1 U20 ( .A1(n44), .A2(n45), .B1(sel[2]), .B2(n46), .ZN(B[0]) );
  INV_X1 U21 ( .A(n46), .ZN(n44) );
  INV_X1 U22 ( .A(AS), .ZN(n45) );
  OAI22_X1 U23 ( .A1(n6), .A2(n38), .B1(n8), .B2(n39), .ZN(B[11]) );
  OAI22_X1 U24 ( .A1(n6), .A2(n21), .B1(n8), .B2(n22), .ZN(B[3]) );
  OAI22_X1 U25 ( .A1(n6), .A2(n13), .B1(n8), .B2(n14), .ZN(B[7]) );
  OAI22_X1 U26 ( .A1(n6), .A2(n28), .B1(n8), .B2(n31), .ZN(B[15]) );
  OAI21_X1 U27 ( .B1(n27), .B2(n28), .A(n29), .ZN(B_17) );
  OR3_X1 U28 ( .A1(A[15]), .A2(n67), .A3(n10), .ZN(n29) );
  AOI21_X1 U29 ( .B1(A[15]), .B2(n67), .A(n30), .ZN(n27) );
  AOI21_X1 U62 ( .B1(n67), .B2(sel[0]), .A(n10), .ZN(AS) );
  NAND2_X1 U63 ( .A1(A[0]), .A2(n30), .ZN(n46) );
  INV_X1 U64 ( .A(n69), .ZN(n68) );
  INV_X1 U65 ( .A(sel[1]), .ZN(n69) );
endmodule


module sum_gen_Nrca4_NB32_0 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_sel_bk_NB4_0 csa_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  carry_sel_bk_NB4_71 csa_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  carry_sel_bk_NB4_70 csa_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  carry_sel_bk_NB4_69 csa_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  carry_sel_bk_NB4_68 csa_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  carry_sel_bk_NB4_67 csa_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  carry_sel_bk_NB4_66 csa_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  carry_sel_bk_NB4_65 csa_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module CSTgen_CW4_NB32_0 ( A, B, Ci, C );
  input [31:0] A;
  input [31:0] B;
  output [7:0] C;
  input Ci;
  wire   g0temp, \matrixProp[0][31] , \matrixProp[0][30] , \matrixProp[0][29] ,
         \matrixProp[0][28] , \matrixProp[0][27] , \matrixProp[0][26] ,
         \matrixProp[0][25] , \matrixProp[0][24] , \matrixProp[0][23] ,
         \matrixProp[0][22] , \matrixProp[0][21] , \matrixProp[0][20] ,
         \matrixProp[0][19] , \matrixProp[0][18] , \matrixProp[0][17] ,
         \matrixProp[0][16] , \matrixProp[0][15] , \matrixProp[0][14] ,
         \matrixProp[0][13] , \matrixProp[0][12] , \matrixProp[0][11] ,
         \matrixProp[0][10] , \matrixProp[0][9] , \matrixProp[0][8] ,
         \matrixProp[0][7] , \matrixProp[0][6] , \matrixProp[0][5] ,
         \matrixProp[0][4] , \matrixProp[0][3] , \matrixProp[0][2] ,
         \matrixProp[0][1] , \matrixProp[0][0] , \matrixProp[1][31] ,
         \matrixProp[1][29] , \matrixProp[1][27] , \matrixProp[1][25] ,
         \matrixProp[1][23] , \matrixProp[1][21] , \matrixProp[1][19] ,
         \matrixProp[1][17] , \matrixProp[1][15] , \matrixProp[1][13] ,
         \matrixProp[1][11] , \matrixProp[1][9] , \matrixProp[1][7] ,
         \matrixProp[1][5] , \matrixProp[1][3] , \matrixProp[2][31] ,
         \matrixProp[2][27] , \matrixProp[2][23] , \matrixProp[2][19] ,
         \matrixProp[2][15] , \matrixProp[2][11] , \matrixProp[2][7] ,
         \matrixProp[3][31] , \matrixProp[3][23] , \matrixProp[3][15] ,
         \matrixProp[4][31] , \matrixProp[4][27] , \matrixGen[0][31] ,
         \matrixGen[0][30] , \matrixGen[0][29] , \matrixGen[0][28] ,
         \matrixGen[0][27] , \matrixGen[0][26] , \matrixGen[0][25] ,
         \matrixGen[0][24] , \matrixGen[0][23] , \matrixGen[0][22] ,
         \matrixGen[0][21] , \matrixGen[0][20] , \matrixGen[0][19] ,
         \matrixGen[0][18] , \matrixGen[0][17] , \matrixGen[0][16] ,
         \matrixGen[0][15] , \matrixGen[0][14] , \matrixGen[0][13] ,
         \matrixGen[0][12] , \matrixGen[0][11] , \matrixGen[0][10] ,
         \matrixGen[0][9] , \matrixGen[0][8] , \matrixGen[0][7] ,
         \matrixGen[0][6] , \matrixGen[0][5] , \matrixGen[0][4] ,
         \matrixGen[0][3] , \matrixGen[0][2] , \matrixGen[0][1] ,
         \matrixGen[1][31] , \matrixGen[1][29] , \matrixGen[1][27] ,
         \matrixGen[1][25] , \matrixGen[1][23] , \matrixGen[1][21] ,
         \matrixGen[1][19] , \matrixGen[1][17] , \matrixGen[1][15] ,
         \matrixGen[1][13] , \matrixGen[1][11] , \matrixGen[1][9] ,
         \matrixGen[1][7] , \matrixGen[1][5] , \matrixGen[1][3] ,
         \matrixGen[1][1] , \matrixGen[2][31] , \matrixGen[2][27] ,
         \matrixGen[2][23] , \matrixGen[2][19] , \matrixGen[2][15] ,
         \matrixGen[2][11] , \matrixGen[2][7] , \matrixGen[3][31] ,
         \matrixGen[3][23] , \matrixGen[3][15] , \matrixGen[4][31] ,
         \matrixGen[4][27] , n7, n4, n2;

  pg_net_0 pg_n0_0 ( .a(A[0]), .b(B[0]), .p(\matrixProp[0][0] ), .g(g0temp) );
  pg_net_287 pg_n_1 ( .a(A[1]), .b(B[1]), .p(\matrixProp[0][1] ), .g(
        \matrixGen[0][1] ) );
  pg_net_286 pg_n_2 ( .a(A[2]), .b(B[2]), .p(\matrixProp[0][2] ), .g(
        \matrixGen[0][2] ) );
  pg_net_285 pg_n_3 ( .a(A[3]), .b(B[3]), .p(\matrixProp[0][3] ), .g(
        \matrixGen[0][3] ) );
  pg_net_284 pg_n_4 ( .a(A[4]), .b(B[4]), .p(\matrixProp[0][4] ), .g(
        \matrixGen[0][4] ) );
  pg_net_283 pg_n_5 ( .a(A[5]), .b(B[5]), .p(\matrixProp[0][5] ), .g(
        \matrixGen[0][5] ) );
  pg_net_282 pg_n_6 ( .a(A[6]), .b(B[6]), .p(\matrixProp[0][6] ), .g(
        \matrixGen[0][6] ) );
  pg_net_281 pg_n_7 ( .a(A[7]), .b(B[7]), .p(\matrixProp[0][7] ), .g(
        \matrixGen[0][7] ) );
  pg_net_280 pg_n_8 ( .a(A[8]), .b(B[8]), .p(\matrixProp[0][8] ), .g(
        \matrixGen[0][8] ) );
  pg_net_279 pg_n_9 ( .a(A[9]), .b(B[9]), .p(\matrixProp[0][9] ), .g(
        \matrixGen[0][9] ) );
  pg_net_278 pg_n_10 ( .a(A[10]), .b(B[10]), .p(\matrixProp[0][10] ), .g(
        \matrixGen[0][10] ) );
  pg_net_277 pg_n_11 ( .a(A[11]), .b(B[11]), .p(\matrixProp[0][11] ), .g(
        \matrixGen[0][11] ) );
  pg_net_276 pg_n_12 ( .a(A[12]), .b(B[12]), .p(\matrixProp[0][12] ), .g(
        \matrixGen[0][12] ) );
  pg_net_275 pg_n_13 ( .a(A[13]), .b(B[13]), .p(\matrixProp[0][13] ), .g(
        \matrixGen[0][13] ) );
  pg_net_274 pg_n_14 ( .a(A[14]), .b(B[14]), .p(\matrixProp[0][14] ), .g(
        \matrixGen[0][14] ) );
  pg_net_273 pg_n_15 ( .a(A[15]), .b(B[15]), .p(\matrixProp[0][15] ), .g(
        \matrixGen[0][15] ) );
  pg_net_272 pg_n_16 ( .a(A[16]), .b(B[16]), .p(\matrixProp[0][16] ), .g(
        \matrixGen[0][16] ) );
  pg_net_271 pg_n_17 ( .a(A[17]), .b(B[17]), .p(\matrixProp[0][17] ), .g(
        \matrixGen[0][17] ) );
  pg_net_270 pg_n_18 ( .a(A[18]), .b(B[18]), .p(\matrixProp[0][18] ), .g(
        \matrixGen[0][18] ) );
  pg_net_269 pg_n_19 ( .a(A[19]), .b(B[19]), .p(\matrixProp[0][19] ), .g(
        \matrixGen[0][19] ) );
  pg_net_268 pg_n_20 ( .a(A[20]), .b(B[20]), .p(\matrixProp[0][20] ), .g(
        \matrixGen[0][20] ) );
  pg_net_267 pg_n_21 ( .a(A[21]), .b(B[21]), .p(\matrixProp[0][21] ), .g(
        \matrixGen[0][21] ) );
  pg_net_266 pg_n_22 ( .a(A[22]), .b(B[22]), .p(\matrixProp[0][22] ), .g(
        \matrixGen[0][22] ) );
  pg_net_265 pg_n_23 ( .a(A[23]), .b(B[23]), .p(\matrixProp[0][23] ), .g(
        \matrixGen[0][23] ) );
  pg_net_264 pg_n_24 ( .a(A[24]), .b(B[24]), .p(\matrixProp[0][24] ), .g(
        \matrixGen[0][24] ) );
  pg_net_263 pg_n_25 ( .a(A[25]), .b(B[25]), .p(\matrixProp[0][25] ), .g(
        \matrixGen[0][25] ) );
  pg_net_262 pg_n_26 ( .a(A[26]), .b(B[26]), .p(\matrixProp[0][26] ), .g(
        \matrixGen[0][26] ) );
  pg_net_261 pg_n_27 ( .a(A[27]), .b(B[27]), .p(\matrixProp[0][27] ), .g(
        \matrixGen[0][27] ) );
  pg_net_260 pg_n_28 ( .a(A[28]), .b(B[28]), .p(\matrixProp[0][28] ), .g(
        \matrixGen[0][28] ) );
  pg_net_259 pg_n_29 ( .a(A[29]), .b(B[29]), .p(\matrixProp[0][29] ), .g(
        \matrixGen[0][29] ) );
  pg_net_258 pg_n_30 ( .a(A[30]), .b(B[30]), .p(\matrixProp[0][30] ), .g(
        \matrixGen[0][30] ) );
  pg_net_257 pg_n_31 ( .a(A[31]), .b(B[31]), .p(\matrixProp[0][31] ), .g(
        \matrixGen[0][31] ) );
  blockPG_0 pg_1_4_0 ( .Gik(\matrixGen[0][3] ), .Gk_1j(\matrixGen[0][2] ), 
        .Pik(\matrixProp[0][3] ), .Pk_1j(\matrixProp[0][2] ), .Pij(
        \matrixProp[1][3] ), .Gij(\matrixGen[1][3] ) );
  G_0 gen_1_4_1 ( .Gik(\matrixGen[0][1] ), .Gk_1j(n4), .Pik(\matrixProp[0][1] ), .Gij(\matrixGen[1][1] ) );
  blockPG_242 pg_1_8_0 ( .Gik(\matrixGen[0][7] ), .Gk_1j(\matrixGen[0][6] ), 
        .Pik(\matrixProp[0][7] ), .Pk_1j(\matrixProp[0][6] ), .Pij(
        \matrixProp[1][7] ), .Gij(\matrixGen[1][7] ) );
  blockPG_241 pg_1_8_1 ( .Gik(\matrixGen[0][5] ), .Gk_1j(\matrixGen[0][4] ), 
        .Pik(\matrixProp[0][5] ), .Pk_1j(\matrixProp[0][4] ), .Pij(
        \matrixProp[1][5] ), .Gij(\matrixGen[1][5] ) );
  blockPG_240 pg_1_12_0 ( .Gik(\matrixGen[0][11] ), .Gk_1j(\matrixGen[0][10] ), 
        .Pik(\matrixProp[0][11] ), .Pk_1j(\matrixProp[0][10] ), .Pij(
        \matrixProp[1][11] ), .Gij(\matrixGen[1][11] ) );
  blockPG_239 pg_1_12_1 ( .Gik(\matrixGen[0][9] ), .Gk_1j(\matrixGen[0][8] ), 
        .Pik(\matrixProp[0][9] ), .Pk_1j(\matrixProp[0][8] ), .Pij(
        \matrixProp[1][9] ), .Gij(\matrixGen[1][9] ) );
  blockPG_238 pg_1_16_0 ( .Gik(\matrixGen[0][15] ), .Gk_1j(\matrixGen[0][14] ), 
        .Pik(\matrixProp[0][15] ), .Pk_1j(\matrixProp[0][14] ), .Pij(
        \matrixProp[1][15] ), .Gij(\matrixGen[1][15] ) );
  blockPG_237 pg_1_16_1 ( .Gik(\matrixGen[0][13] ), .Gk_1j(\matrixGen[0][12] ), 
        .Pik(\matrixProp[0][13] ), .Pk_1j(\matrixProp[0][12] ), .Pij(
        \matrixProp[1][13] ), .Gij(\matrixGen[1][13] ) );
  blockPG_236 pg_1_20_0 ( .Gik(\matrixGen[0][19] ), .Gk_1j(\matrixGen[0][18] ), 
        .Pik(\matrixProp[0][19] ), .Pk_1j(\matrixProp[0][18] ), .Pij(
        \matrixProp[1][19] ), .Gij(\matrixGen[1][19] ) );
  blockPG_235 pg_1_20_1 ( .Gik(\matrixGen[0][17] ), .Gk_1j(\matrixGen[0][16] ), 
        .Pik(\matrixProp[0][17] ), .Pk_1j(\matrixProp[0][16] ), .Pij(
        \matrixProp[1][17] ), .Gij(\matrixGen[1][17] ) );
  blockPG_234 pg_1_24_0 ( .Gik(\matrixGen[0][23] ), .Gk_1j(\matrixGen[0][22] ), 
        .Pik(\matrixProp[0][23] ), .Pk_1j(\matrixProp[0][22] ), .Pij(
        \matrixProp[1][23] ), .Gij(\matrixGen[1][23] ) );
  blockPG_233 pg_1_24_1 ( .Gik(\matrixGen[0][21] ), .Gk_1j(\matrixGen[0][20] ), 
        .Pik(\matrixProp[0][21] ), .Pk_1j(\matrixProp[0][20] ), .Pij(
        \matrixProp[1][21] ), .Gij(\matrixGen[1][21] ) );
  blockPG_232 pg_1_28_0 ( .Gik(\matrixGen[0][27] ), .Gk_1j(\matrixGen[0][26] ), 
        .Pik(\matrixProp[0][27] ), .Pk_1j(\matrixProp[0][26] ), .Pij(
        \matrixProp[1][27] ), .Gij(\matrixGen[1][27] ) );
  blockPG_231 pg_1_28_1 ( .Gik(\matrixGen[0][25] ), .Gk_1j(\matrixGen[0][24] ), 
        .Pik(\matrixProp[0][25] ), .Pk_1j(\matrixProp[0][24] ), .Pij(
        \matrixProp[1][25] ), .Gij(\matrixGen[1][25] ) );
  blockPG_230 pg_1_32_0 ( .Gik(\matrixGen[0][31] ), .Gk_1j(\matrixGen[0][30] ), 
        .Pik(\matrixProp[0][31] ), .Pk_1j(\matrixProp[0][30] ), .Pij(
        \matrixProp[1][31] ), .Gij(\matrixGen[1][31] ) );
  blockPG_229 pg_1_32_1 ( .Gik(\matrixGen[0][29] ), .Gk_1j(\matrixGen[0][28] ), 
        .Pik(\matrixProp[0][29] ), .Pk_1j(\matrixProp[0][28] ), .Pij(
        \matrixProp[1][29] ), .Gij(\matrixGen[1][29] ) );
  G_80 gen_2_4_0 ( .Gik(\matrixGen[1][3] ), .Gk_1j(\matrixGen[1][1] ), .Pik(
        \matrixProp[1][3] ), .Gij(n7) );
  blockPG_228 pg_2_8_0 ( .Gik(\matrixGen[1][7] ), .Gk_1j(\matrixGen[1][5] ), 
        .Pik(\matrixProp[1][7] ), .Pk_1j(\matrixProp[1][5] ), .Pij(
        \matrixProp[2][7] ), .Gij(\matrixGen[2][7] ) );
  blockPG_227 pg_2_12_0 ( .Gik(\matrixGen[1][11] ), .Gk_1j(\matrixGen[1][9] ), 
        .Pik(\matrixProp[1][11] ), .Pk_1j(\matrixProp[1][9] ), .Pij(
        \matrixProp[2][11] ), .Gij(\matrixGen[2][11] ) );
  blockPG_226 pg_2_16_0 ( .Gik(\matrixGen[1][15] ), .Gk_1j(\matrixGen[1][13] ), 
        .Pik(\matrixProp[1][15] ), .Pk_1j(\matrixProp[1][13] ), .Pij(
        \matrixProp[2][15] ), .Gij(\matrixGen[2][15] ) );
  blockPG_225 pg_2_20_0 ( .Gik(\matrixGen[1][19] ), .Gk_1j(\matrixGen[1][17] ), 
        .Pik(\matrixProp[1][19] ), .Pk_1j(\matrixProp[1][17] ), .Pij(
        \matrixProp[2][19] ), .Gij(\matrixGen[2][19] ) );
  blockPG_224 pg_2_24_0 ( .Gik(\matrixGen[1][23] ), .Gk_1j(\matrixGen[1][21] ), 
        .Pik(\matrixProp[1][23] ), .Pk_1j(\matrixProp[1][21] ), .Pij(
        \matrixProp[2][23] ), .Gij(\matrixGen[2][23] ) );
  blockPG_223 pg_2_28_0 ( .Gik(\matrixGen[1][27] ), .Gk_1j(\matrixGen[1][25] ), 
        .Pik(\matrixProp[1][27] ), .Pk_1j(\matrixProp[1][25] ), .Pij(
        \matrixProp[2][27] ), .Gij(\matrixGen[2][27] ) );
  blockPG_222 pg_2_32_0 ( .Gik(\matrixGen[1][31] ), .Gk_1j(\matrixGen[1][29] ), 
        .Pik(\matrixProp[1][31] ), .Pk_1j(\matrixProp[1][29] ), .Pij(
        \matrixProp[2][31] ), .Gij(\matrixGen[2][31] ) );
  G_79 gen2_3_8_1 ( .Gik(\matrixGen[2][7] ), .Gk_1j(n7), .Pik(
        \matrixProp[2][7] ), .Gij(C[1]) );
  blockPG_221 pg1_3_16_1 ( .Gik(\matrixGen[2][15] ), .Gk_1j(\matrixGen[2][11] ), .Pik(\matrixProp[2][15] ), .Pk_1j(\matrixProp[2][11] ), .Pij(
        \matrixProp[3][15] ), .Gij(\matrixGen[3][15] ) );
  blockPG_220 pg1_3_24_1 ( .Gik(\matrixGen[2][23] ), .Gk_1j(\matrixGen[2][19] ), .Pik(\matrixProp[2][23] ), .Pk_1j(\matrixProp[2][19] ), .Pij(
        \matrixProp[3][23] ), .Gij(\matrixGen[3][23] ) );
  blockPG_219 pg1_3_32_1 ( .Gik(\matrixGen[2][31] ), .Gk_1j(\matrixGen[2][27] ), .Pik(\matrixProp[2][31] ), .Pk_1j(\matrixProp[2][27] ), .Pij(
        \matrixProp[3][31] ), .Gij(\matrixGen[3][31] ) );
  G_78 gen2_4_16_1 ( .Gik(\matrixGen[3][15] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[3][15] ), .Gij(C[3]) );
  G_77 gen2_4_16_2 ( .Gik(\matrixGen[2][11] ), .Gk_1j(C[1]), .Pik(
        \matrixProp[2][11] ), .Gij(C[2]) );
  blockPG_218 pg1_4_32_1 ( .Gik(\matrixGen[3][31] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[3][31] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][31] ), .Gij(\matrixGen[4][31] ) );
  blockPG_217 pg1_4_32_2 ( .Gik(\matrixGen[2][27] ), .Gk_1j(\matrixGen[3][23] ), .Pik(\matrixProp[2][27] ), .Pk_1j(\matrixProp[3][23] ), .Pij(
        \matrixProp[4][27] ), .Gij(\matrixGen[4][27] ) );
  G_76 gen2_5_32_1 ( .Gik(\matrixGen[4][31] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][31] ), .Gij(C[7]) );
  G_75 gen2_5_32_2 ( .Gik(\matrixGen[4][27] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[4][27] ), .Gij(C[6]) );
  G_74 gen2_5_32_3 ( .Gik(\matrixGen[3][23] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[3][23] ), .Gij(C[5]) );
  G_73 gen2_5_32_4 ( .Gik(\matrixGen[2][19] ), .Gk_1j(C[3]), .Pik(
        \matrixProp[2][19] ), .Gij(C[4]) );
  CLKBUF_X1 U1 ( .A(n7), .Z(C[0]) );
  INV_X1 U2 ( .A(n2), .ZN(n4) );
  AOI21_X1 U3 ( .B1(\matrixProp[0][0] ), .B2(Ci), .A(g0temp), .ZN(n2) );
endmodule


module BP_NB32_BP_LEN4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n35,
         n36, n37, n38, n39, n40, n41, n42, n55, n56, n57, n58, n59, n60, n128,
         n129, n145, n149, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n170, n171, n172,
         n173, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318;

  BUF_X2 U2 ( .A(B[31]), .Z(n225) );
  BUF_X2 U3 ( .A(B[31]), .Z(n224) );
  AND3_X1 U4 ( .A1(n311), .A2(n267), .A3(n264), .ZN(n214) );
  XOR2_X1 U5 ( .A(n221), .B(n273), .Z(SUM[29]) );
  NAND2_X1 U6 ( .A1(n183), .A2(n184), .ZN(n181) );
  NAND2_X1 U7 ( .A1(n4), .A2(n12), .ZN(n184) );
  INV_X1 U8 ( .A(n27), .ZN(n24) );
  OAI21_X1 U9 ( .B1(n176), .B2(n157), .A(n159), .ZN(n173) );
  INV_X1 U10 ( .A(n177), .ZN(n176) );
  OAI21_X1 U11 ( .B1(n193), .B2(n200), .A(n10), .ZN(n198) );
  INV_X1 U12 ( .A(n8), .ZN(n200) );
  OAI21_X1 U13 ( .B1(n179), .B2(n180), .A(n158), .ZN(n177) );
  INV_X1 U14 ( .A(n161), .ZN(n179) );
  INV_X1 U15 ( .A(n181), .ZN(n180) );
  OAI21_X1 U16 ( .B1(n29), .B2(n207), .A(n30), .ZN(n27) );
  INV_X1 U17 ( .A(n31), .ZN(n29) );
  INV_X1 U18 ( .A(n41), .ZN(n208) );
  INV_X1 U19 ( .A(n39), .ZN(n212) );
  NAND2_X1 U20 ( .A1(n12), .A2(n14), .ZN(n201) );
  XNOR2_X1 U21 ( .A(n215), .B(n243), .ZN(SUM[27]) );
  NAND2_X1 U22 ( .A1(n232), .A2(n233), .ZN(n215) );
  OAI21_X1 U23 ( .B1(n196), .B2(n197), .A(n192), .ZN(n195) );
  INV_X1 U24 ( .A(n186), .ZN(n197) );
  INV_X1 U25 ( .A(n198), .ZN(n196) );
  OAI21_X1 U26 ( .B1(n37), .B2(n38), .A(n39), .ZN(n36) );
  INV_X1 U27 ( .A(n60), .ZN(n38) );
  INV_X1 U28 ( .A(n40), .ZN(n37) );
  AND2_X1 U29 ( .A1(n304), .A2(n232), .ZN(n216) );
  OAI21_X1 U30 ( .B1(n187), .B2(n188), .A(n189), .ZN(n164) );
  INV_X1 U31 ( .A(n185), .ZN(n188) );
  INV_X1 U32 ( .A(n192), .ZN(n191) );
  OAI21_X1 U33 ( .B1(n157), .B2(n158), .A(n159), .ZN(n154) );
  AOI21_X1 U34 ( .B1(n153), .B2(n154), .A(n155), .ZN(n149) );
  NAND2_X1 U35 ( .A1(n17), .A2(n18), .ZN(n16) );
  NAND2_X1 U36 ( .A1(n19), .A2(n20), .ZN(n17) );
  NAND2_X1 U37 ( .A1(n172), .A2(n156), .ZN(n171) );
  NAND2_X1 U38 ( .A1(n153), .A2(n173), .ZN(n172) );
  NAND2_X1 U39 ( .A1(n19), .A2(n18), .ZN(n23) );
  NAND2_X1 U40 ( .A1(n156), .A2(n153), .ZN(n175) );
  INV_X1 U41 ( .A(n162), .ZN(n157) );
  NAND2_X1 U42 ( .A1(n13), .A2(n14), .ZN(n11) );
  NAND2_X1 U43 ( .A1(n9), .A2(n10), .ZN(n7) );
  INV_X1 U44 ( .A(n21), .ZN(n204) );
  NAND2_X1 U45 ( .A1(n192), .A2(n186), .ZN(n199) );
  NAND2_X1 U46 ( .A1(n159), .A2(n162), .ZN(n178) );
  NAND2_X1 U47 ( .A1(n158), .A2(n161), .ZN(n182) );
  NAND2_X1 U48 ( .A1(n41), .A2(n42), .ZN(n35) );
  NAND2_X1 U49 ( .A1(n21), .A2(n22), .ZN(n15) );
  NAND2_X1 U50 ( .A1(n30), .A2(n31), .ZN(n33) );
  NAND2_X1 U51 ( .A1(n60), .A2(n39), .ZN(n55) );
  NAND2_X1 U52 ( .A1(n189), .A2(n185), .ZN(n194) );
  AND4_X1 U53 ( .A1(n185), .A2(n186), .A3(n9), .A4(n14), .ZN(n4) );
  INV_X1 U54 ( .A(n9), .ZN(n193) );
  BUF_X1 U55 ( .A(B[31]), .Z(n226) );
  INV_X1 U56 ( .A(n156), .ZN(n155) );
  INV_X1 U57 ( .A(n18), .ZN(n206) );
  AND3_X1 U58 ( .A1(n153), .A2(n161), .A3(n162), .ZN(n217) );
  XNOR2_X1 U59 ( .A(n7), .B(n8), .ZN(SUM[9]) );
  NAND2_X1 U60 ( .A1(B[6]), .A2(A[6]), .ZN(n18) );
  NAND2_X1 U61 ( .A1(B[14]), .A2(A[14]), .ZN(n156) );
  NAND2_X1 U62 ( .A1(B[10]), .A2(A[10]), .ZN(n192) );
  NAND2_X1 U63 ( .A1(B[12]), .A2(A[12]), .ZN(n158) );
  NAND2_X1 U64 ( .A1(B[13]), .A2(A[13]), .ZN(n159) );
  NAND2_X1 U65 ( .A1(B[9]), .A2(A[9]), .ZN(n10) );
  NAND2_X1 U66 ( .A1(B[4]), .A2(A[4]), .ZN(n30) );
  OR2_X1 U67 ( .A1(B[10]), .A2(A[10]), .ZN(n186) );
  NAND2_X1 U68 ( .A1(B[11]), .A2(A[11]), .ZN(n189) );
  XNOR2_X1 U69 ( .A(n170), .B(n171), .ZN(SUM[15]) );
  NAND2_X1 U70 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U71 ( .A1(B[7]), .A2(A[7]), .ZN(n22) );
  NAND2_X1 U72 ( .A1(B[3]), .A2(A[3]), .ZN(n42) );
  OR2_X1 U73 ( .A1(B[8]), .A2(A[8]), .ZN(n14) );
  OR2_X1 U74 ( .A1(B[6]), .A2(A[6]), .ZN(n19) );
  OR2_X1 U75 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OR2_X1 U76 ( .A1(B[11]), .A2(A[11]), .ZN(n185) );
  OR2_X1 U77 ( .A1(B[4]), .A2(A[4]), .ZN(n31) );
  OR2_X1 U78 ( .A1(B[7]), .A2(A[7]), .ZN(n21) );
  NAND2_X1 U79 ( .A1(n56), .A2(n57), .ZN(n40) );
  OR2_X1 U80 ( .A1(B[3]), .A2(A[3]), .ZN(n41) );
  OR2_X1 U81 ( .A1(B[5]), .A2(A[5]), .ZN(n32) );
  XNOR2_X1 U82 ( .A(n194), .B(n195), .ZN(SUM[11]) );
  XNOR2_X1 U83 ( .A(n199), .B(n198), .ZN(SUM[10]) );
  XNOR2_X1 U84 ( .A(n35), .B(n36), .ZN(SUM[3]) );
  XNOR2_X1 U85 ( .A(n33), .B(n167), .ZN(SUM[4]) );
  XNOR2_X1 U86 ( .A(n23), .B(n20), .ZN(SUM[6]) );
  XNOR2_X1 U87 ( .A(n15), .B(n16), .ZN(SUM[7]) );
  XNOR2_X1 U88 ( .A(n175), .B(n173), .ZN(SUM[14]) );
  XNOR2_X1 U89 ( .A(n178), .B(n177), .ZN(SUM[13]) );
  XNOR2_X1 U90 ( .A(n55), .B(n40), .ZN(SUM[2]) );
  XNOR2_X1 U91 ( .A(n28), .B(n27), .ZN(SUM[5]) );
  XNOR2_X1 U92 ( .A(n182), .B(n181), .ZN(SUM[12]) );
  XNOR2_X1 U93 ( .A(n11), .B(n12), .ZN(SUM[8]) );
  INV_X1 U94 ( .A(n220), .ZN(n58) );
  XNOR2_X1 U95 ( .A(n128), .B(n59), .ZN(SUM[1]) );
  OR2_X1 U96 ( .A1(B[0]), .A2(A[0]), .ZN(n209) );
  OAI21_X1 U97 ( .B1(n24), .B2(n25), .A(n26), .ZN(n20) );
  NAND2_X1 U98 ( .A1(n287), .A2(n214), .ZN(n313) );
  NAND2_X1 U99 ( .A1(n32), .A2(n26), .ZN(n28) );
  NAND2_X1 U100 ( .A1(n299), .A2(n217), .ZN(n308) );
  OR2_X1 U101 ( .A1(B[13]), .A2(A[13]), .ZN(n162) );
  OR2_X1 U102 ( .A1(B[12]), .A2(A[12]), .ZN(n161) );
  OR2_X1 U103 ( .A1(B[14]), .A2(A[14]), .ZN(n153) );
  NAND2_X1 U104 ( .A1(B[5]), .A2(A[5]), .ZN(n26) );
  INV_X1 U105 ( .A(n261), .ZN(n218) );
  NAND2_X1 U106 ( .A1(n281), .A2(n219), .ZN(n234) );
  NOR2_X1 U107 ( .A1(n235), .A2(n218), .ZN(n219) );
  AND2_X1 U108 ( .A1(n129), .A2(n209), .ZN(SUM[0]) );
  AOI21_X1 U109 ( .B1(n186), .B2(n190), .A(n191), .ZN(n187) );
  NAND2_X1 U110 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  OAI21_X1 U111 ( .B1(n193), .B2(n13), .A(n10), .ZN(n190) );
  NAND2_X1 U112 ( .A1(n201), .A2(n13), .ZN(n8) );
  OAI21_X1 U113 ( .B1(n207), .B2(n168), .A(n165), .ZN(n12) );
  INV_X1 U114 ( .A(n168), .ZN(n160) );
  NAND2_X1 U115 ( .A1(B[0]), .A2(A[0]), .ZN(n129) );
  INV_X1 U116 ( .A(n129), .ZN(n59) );
  INV_X1 U117 ( .A(n164), .ZN(n183) );
  NOR2_X1 U118 ( .A1(B[1]), .A2(A[1]), .ZN(n220) );
  NAND4_X1 U119 ( .A1(n31), .A2(n32), .A3(n19), .A4(n21), .ZN(n168) );
  INV_X1 U120 ( .A(n32), .ZN(n25) );
  NAND2_X1 U121 ( .A1(n58), .A2(n57), .ZN(n128) );
  NAND2_X1 U122 ( .A1(n58), .A2(n59), .ZN(n56) );
  NAND2_X1 U123 ( .A1(n315), .A2(n216), .ZN(n275) );
  AOI21_X1 U124 ( .B1(n306), .B2(n275), .A(n242), .ZN(n221) );
  OR2_X1 U125 ( .A1(B[2]), .A2(A[2]), .ZN(n60) );
  NOR2_X1 U126 ( .A1(n286), .A2(n270), .ZN(n222) );
  OAI21_X1 U127 ( .B1(n221), .B2(n292), .A(n293), .ZN(n223) );
  NAND2_X1 U128 ( .A1(B[1]), .A2(A[1]), .ZN(n57) );
  OAI21_X1 U129 ( .B1(n25), .B2(n30), .A(n26), .ZN(n205) );
  INV_X1 U130 ( .A(n202), .ZN(n165) );
  INV_X1 U131 ( .A(n167), .ZN(n207) );
  NAND2_X1 U132 ( .A1(n160), .A2(n167), .ZN(n166) );
  OAI21_X1 U133 ( .B1(n210), .B2(n208), .A(n42), .ZN(n167) );
  OAI21_X1 U134 ( .B1(n220), .B2(n129), .A(n57), .ZN(n211) );
  AOI21_X1 U135 ( .B1(n4), .B2(n163), .A(n164), .ZN(n145) );
  NAND2_X1 U136 ( .A1(n165), .A2(n166), .ZN(n163) );
  AOI21_X1 U137 ( .B1(n211), .B2(n60), .A(n212), .ZN(n210) );
  OAI21_X1 U138 ( .B1(n203), .B2(n204), .A(n22), .ZN(n202) );
  AOI21_X1 U139 ( .B1(n205), .B2(n19), .A(n206), .ZN(n203) );
  NAND2_X1 U140 ( .A1(n227), .A2(n228), .ZN(n170) );
  NOR2_X1 U141 ( .A1(n230), .A2(n231), .ZN(n229) );
  NOR2_X1 U142 ( .A1(n238), .A2(n239), .ZN(n237) );
  NOR2_X1 U143 ( .A1(n241), .A2(n242), .ZN(n240) );
  AOI21_X1 U144 ( .B1(n244), .B2(n245), .A(n246), .ZN(n243) );
  AND2_X1 U145 ( .A1(n248), .A2(n249), .ZN(n247) );
  NOR2_X1 U146 ( .A1(n251), .A2(n252), .ZN(n250) );
  AOI21_X1 U147 ( .B1(n254), .B2(n255), .A(n256), .ZN(n253) );
  NOR2_X1 U148 ( .A1(n258), .A2(n259), .ZN(n257) );
  AND2_X1 U149 ( .A1(n261), .A2(n262), .ZN(n260) );
  AND2_X1 U150 ( .A1(n264), .A2(n265), .ZN(n263) );
  AND2_X1 U151 ( .A1(n267), .A2(n268), .ZN(n266) );
  NOR2_X1 U152 ( .A1(n270), .A2(n271), .ZN(n269) );
  XOR2_X1 U153 ( .A(n223), .B(n237), .Z(SUM[30]) );
  XOR2_X1 U154 ( .A(n275), .B(n240), .Z(SUM[28]) );
  XOR2_X1 U155 ( .A(n276), .B(n244), .Z(SUM[26]) );
  XNOR2_X1 U156 ( .A(n277), .B(n247), .ZN(SUM[25]) );
  XOR2_X1 U157 ( .A(n278), .B(n250), .Z(SUM[24]) );
  XOR2_X1 U158 ( .A(n279), .B(n254), .Z(SUM[22]) );
  XOR2_X1 U159 ( .A(n280), .B(n257), .Z(SUM[21]) );
  XOR2_X1 U160 ( .A(n281), .B(n260), .Z(SUM[20]) );
  XOR2_X1 U161 ( .A(n282), .B(n263), .Z(SUM[19]) );
  XOR2_X1 U162 ( .A(n283), .B(n284), .Z(SUM[18]) );
  XNOR2_X1 U163 ( .A(n285), .B(n266), .ZN(SUM[17]) );
  XNOR2_X1 U164 ( .A(n286), .B(n269), .ZN(SUM[16]) );
  NOR2_X1 U165 ( .A1(n286), .A2(n270), .ZN(n287) );
  OR3_X1 U166 ( .A1(n258), .A2(n256), .A3(n230), .ZN(n235) );
  NAND2_X1 U167 ( .A1(n281), .A2(n261), .ZN(n236) );
  AND4_X1 U168 ( .A1(n289), .A2(n290), .A3(n255), .A4(n262), .ZN(n288) );
  AOI21_X1 U169 ( .B1(n234), .B2(n288), .A(n251), .ZN(n291) );
  OAI21_X1 U170 ( .B1(n274), .B2(n292), .A(n293), .ZN(n272) );
  OAI21_X1 U171 ( .B1(n295), .B2(n277), .A(n249), .ZN(n294) );
  AOI21_X1 U172 ( .B1(n296), .B2(n280), .A(n259), .ZN(n254) );
  XOR2_X1 U173 ( .A(n297), .B(n298), .Z(SUM[31]) );
  XOR2_X1 U174 ( .A(n229), .B(n253), .Z(SUM[23]) );
  NOR2_X1 U175 ( .A1(n145), .A2(n300), .ZN(n299) );
  AND3_X1 U176 ( .A1(n268), .A2(n302), .A3(n303), .ZN(n301) );
  AND3_X1 U177 ( .A1(n249), .A2(n305), .A3(n245), .ZN(n304) );
  AOI21_X1 U178 ( .B1(n306), .B2(n275), .A(n242), .ZN(n274) );
  NAND2_X1 U179 ( .A1(n225), .A2(A[15]), .ZN(n227) );
  NOR2_X1 U180 ( .A1(n224), .A2(A[15]), .ZN(n300) );
  INV_X1 U181 ( .A(n300), .ZN(n228) );
  AND2_X1 U182 ( .A1(A[28]), .A2(n226), .ZN(n242) );
  NAND2_X1 U183 ( .A1(A[24]), .A2(n225), .ZN(n305) );
  INV_X1 U184 ( .A(n305), .ZN(n252) );
  NAND2_X1 U185 ( .A1(A[26]), .A2(n225), .ZN(n245) );
  NAND2_X1 U186 ( .A1(A[25]), .A2(n225), .ZN(n249) );
  NAND2_X1 U187 ( .A1(A[27]), .A2(n225), .ZN(n232) );
  NOR2_X1 U188 ( .A1(n224), .A2(A[26]), .ZN(n246) );
  INV_X1 U189 ( .A(n246), .ZN(n307) );
  NOR2_X1 U190 ( .A1(n224), .A2(A[25]), .ZN(n295) );
  OR2_X1 U191 ( .A1(n226), .A2(A[27]), .ZN(n233) );
  NOR2_X1 U192 ( .A1(n224), .A2(A[24]), .ZN(n251) );
  OAI211_X1 U193 ( .C1(n149), .C2(n300), .A(n227), .B(n308), .ZN(n309) );
  NOR2_X1 U194 ( .A1(n224), .A2(A[16]), .ZN(n270) );
  NOR2_X1 U195 ( .A1(n224), .A2(A[18]), .ZN(n310) );
  INV_X1 U196 ( .A(n310), .ZN(n311) );
  NOR2_X1 U197 ( .A1(n224), .A2(A[17]), .ZN(n312) );
  OR2_X1 U198 ( .A1(n226), .A2(A[19]), .ZN(n264) );
  NAND2_X1 U199 ( .A1(A[16]), .A2(n225), .ZN(n302) );
  INV_X1 U200 ( .A(n302), .ZN(n271) );
  NAND2_X1 U201 ( .A1(A[18]), .A2(n225), .ZN(n303) );
  NAND2_X1 U202 ( .A1(A[17]), .A2(n225), .ZN(n268) );
  NAND2_X1 U203 ( .A1(A[19]), .A2(n225), .ZN(n265) );
  NAND3_X1 U204 ( .A1(n313), .A2(n265), .A3(n301), .ZN(n281) );
  OR2_X1 U205 ( .A1(n226), .A2(A[20]), .ZN(n261) );
  NOR2_X1 U206 ( .A1(n224), .A2(A[22]), .ZN(n256) );
  INV_X1 U207 ( .A(n256), .ZN(n314) );
  NOR2_X1 U208 ( .A1(n224), .A2(A[21]), .ZN(n258) );
  NOR2_X1 U209 ( .A1(n224), .A2(A[23]), .ZN(n230) );
  NAND2_X1 U210 ( .A1(A[20]), .A2(n225), .ZN(n262) );
  NAND2_X1 U211 ( .A1(A[22]), .A2(n225), .ZN(n255) );
  NAND2_X1 U212 ( .A1(A[21]), .A2(n225), .ZN(n290) );
  INV_X1 U213 ( .A(n290), .ZN(n259) );
  NAND2_X1 U214 ( .A1(A[23]), .A2(n225), .ZN(n289) );
  INV_X1 U215 ( .A(n289), .ZN(n231) );
  NAND4_X1 U216 ( .A1(n291), .A2(n233), .A3(n248), .A4(n307), .ZN(n315) );
  NOR2_X1 U217 ( .A1(n224), .A2(A[28]), .ZN(n241) );
  NAND2_X1 U218 ( .A1(A[29]), .A2(n225), .ZN(n293) );
  NOR2_X1 U219 ( .A1(n224), .A2(A[29]), .ZN(n292) );
  INV_X1 U220 ( .A(n292), .ZN(n316) );
  NOR2_X1 U221 ( .A1(n224), .A2(A[30]), .ZN(n239) );
  INV_X1 U222 ( .A(n239), .ZN(n317) );
  AND2_X1 U223 ( .A1(A[30]), .A2(n226), .ZN(n238) );
  OAI21_X1 U224 ( .B1(n238), .B2(n272), .A(n317), .ZN(n297) );
  NAND2_X1 U225 ( .A1(n293), .A2(n316), .ZN(n273) );
  NOR2_X1 U226 ( .A1(n252), .A2(n291), .ZN(n277) );
  NAND2_X1 U227 ( .A1(n307), .A2(n245), .ZN(n276) );
  OAI21_X1 U228 ( .B1(n235), .B2(n236), .A(n288), .ZN(n278) );
  NAND2_X1 U229 ( .A1(n262), .A2(n236), .ZN(n280) );
  NAND2_X1 U230 ( .A1(n314), .A2(n255), .ZN(n279) );
  NOR2_X1 U231 ( .A1(n271), .A2(n222), .ZN(n285) );
  OAI21_X1 U232 ( .B1(n312), .B2(n285), .A(n268), .ZN(n318) );
  OAI21_X1 U233 ( .B1(n284), .B2(n310), .A(n303), .ZN(n282) );
  NAND2_X1 U234 ( .A1(n303), .A2(n311), .ZN(n283) );
  XNOR2_X1 U235 ( .A(n224), .B(A[31]), .ZN(n298) );
  INV_X1 U236 ( .A(n309), .ZN(n286) );
  INV_X1 U237 ( .A(n241), .ZN(n306) );
  INV_X1 U238 ( .A(n295), .ZN(n248) );
  INV_X1 U239 ( .A(n258), .ZN(n296) );
  INV_X1 U240 ( .A(n312), .ZN(n267) );
  INV_X1 U241 ( .A(n294), .ZN(n244) );
  INV_X1 U242 ( .A(n318), .ZN(n284) );
endmodule


module BP_NB32_BP_LEN4_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
  NOR4_X1 U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(EQ) );
  NAND4_X1 U2 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n18), .A2(n19), .ZN(n2) );
  NAND4_X1 U4 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n1) );
  NOR4_X1 U5 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  NOR4_X1 U6 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  NOR4_X1 U7 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  NOR4_X1 U8 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  NOR4_X1 U9 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  NOR4_X1 U10 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  OAI22_X1 U11 ( .A1(n13), .A2(n14), .B1(B[1]), .B2(n13), .ZN(n12) );
  INV_X1 U12 ( .A(A[1]), .ZN(n14) );
  AND2_X1 U13 ( .A1(B[0]), .A2(n15), .ZN(n13) );
  NOR2_X1 U14 ( .A1(n15), .A2(B[0]), .ZN(n16) );
  XNOR2_X1 U15 ( .A(B[3]), .B(A[3]), .ZN(n8) );
  XNOR2_X1 U16 ( .A(B[6]), .B(A[6]), .ZN(n5) );
  INV_X1 U17 ( .A(B[1]), .ZN(n17) );
  NAND4_X1 U18 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  XNOR2_X1 U23 ( .A(B[2]), .B(A[2]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(A[1]), .A2(n16), .B1(n16), .B2(n17), .ZN(n11) );
  XNOR2_X1 U29 ( .A(B[31]), .B(A[31]), .ZN(n10) );
  XNOR2_X1 U34 ( .A(B[4]), .B(A[4]), .ZN(n7) );
  XNOR2_X1 U39 ( .A(B[5]), .B(A[5]), .ZN(n6) );
  INV_X1 U44 ( .A(A[0]), .ZN(n15) );
endmodule


module BP_NB32_BP_LEN4_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n29, n30, n31, n32, n33, n34,
         n35, n36, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;

  XOR2_X1 U20 ( .A(B[10]), .B(A[10]), .Z(n24) );
  XOR2_X1 U21 ( .A(B[9]), .B(A[9]), .Z(n23) );
  XOR2_X1 U22 ( .A(B[8]), .B(A[8]), .Z(n22) );
  XOR2_X1 U23 ( .A(B[7]), .B(A[7]), .Z(n21) );
  XOR2_X1 U31 ( .A(B[18]), .B(A[18]), .Z(n36) );
  XOR2_X1 U32 ( .A(B[17]), .B(A[17]), .Z(n35) );
  XOR2_X1 U33 ( .A(B[16]), .B(A[16]), .Z(n34) );
  XOR2_X1 U34 ( .A(B[15]), .B(A[15]), .Z(n33) );
  INV_X1 U1 ( .A(B[1]), .ZN(n18) );
  NOR2_X1 U2 ( .A1(n16), .A2(B[0]), .ZN(n17) );
  OR3_X1 U3 ( .A1(n3), .A2(n4), .A3(n5), .ZN(n1) );
  NAND4_X1 U4 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  AND2_X1 U5 ( .A1(B[0]), .A2(n16), .ZN(n14) );
  NOR4_X1 U6 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .ZN(n32) );
  XNOR2_X1 U7 ( .A(B[6]), .B(A[6]), .ZN(n6) );
  XNOR2_X1 U8 ( .A(B[4]), .B(A[4]), .ZN(n8) );
  XNOR2_X1 U9 ( .A(B[3]), .B(A[3]), .ZN(n9) );
  XNOR2_X1 U10 ( .A(B[5]), .B(A[5]), .ZN(n7) );
  NAND4_X1 U11 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(n4) );
  OAI22_X1 U12 ( .A1(n14), .A2(n15), .B1(B[1]), .B2(n14), .ZN(n13) );
  XNOR2_X1 U13 ( .A(B[2]), .B(A[2]), .ZN(n10) );
  OAI22_X1 U14 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n18), .ZN(n12) );
  NOR4_X1 U15 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n20) );
  AND4_X1 U16 ( .A1(n59), .A2(n58), .A3(n57), .A4(n60), .ZN(n31) );
  INV_X1 U17 ( .A(A[0]), .ZN(n16) );
  INV_X1 U18 ( .A(A[1]), .ZN(n15) );
  AND4_X1 U19 ( .A1(n49), .A2(n50), .A3(n51), .A4(n52), .ZN(n19) );
  XNOR2_X1 U24 ( .A(B[11]), .B(A[11]), .ZN(n49) );
  XNOR2_X1 U25 ( .A(B[12]), .B(A[12]), .ZN(n50) );
  XNOR2_X1 U26 ( .A(B[13]), .B(A[13]), .ZN(n51) );
  XNOR2_X1 U27 ( .A(B[14]), .B(A[14]), .ZN(n52) );
  XNOR2_X1 U28 ( .A(B[31]), .B(A[31]), .ZN(n11) );
  AND4_X1 U29 ( .A1(n53), .A2(n54), .A3(n55), .A4(n56), .ZN(n29) );
  XNOR2_X1 U30 ( .A(B[27]), .B(A[27]), .ZN(n53) );
  XNOR2_X1 U35 ( .A(B[28]), .B(A[28]), .ZN(n54) );
  XNOR2_X1 U36 ( .A(B[29]), .B(A[29]), .ZN(n55) );
  XNOR2_X1 U37 ( .A(B[30]), .B(A[30]), .ZN(n56) );
  XNOR2_X1 U38 ( .A(B[19]), .B(A[19]), .ZN(n57) );
  XNOR2_X1 U39 ( .A(B[20]), .B(A[20]), .ZN(n58) );
  XNOR2_X1 U40 ( .A(B[21]), .B(A[21]), .ZN(n59) );
  XNOR2_X1 U41 ( .A(B[22]), .B(A[22]), .ZN(n60) );
  AND4_X1 U42 ( .A1(n61), .A2(n62), .A3(n63), .A4(n64), .ZN(n30) );
  XNOR2_X1 U43 ( .A(B[23]), .B(A[23]), .ZN(n61) );
  XNOR2_X1 U44 ( .A(B[24]), .B(A[24]), .ZN(n62) );
  XNOR2_X1 U45 ( .A(B[25]), .B(A[25]), .ZN(n63) );
  XNOR2_X1 U46 ( .A(B[26]), .B(A[26]), .ZN(n64) );
  NAND2_X1 U47 ( .A1(n19), .A2(n20), .ZN(n3) );
  NOR2_X1 U48 ( .A1(n2), .A2(n1), .ZN(EQ) );
  NAND4_X1 U49 ( .A1(n29), .A2(n30), .A3(n31), .A4(n32), .ZN(n2) );
endmodule


module FD_NB5_1 ( CK, RESET, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
endmodule


module EXECUTION_UNIT_NB32_LS5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , n1;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X1 U3 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  XOR2_X1 U5 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  XOR2_X1 U7 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  XOR2_X1 U9 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  XOR2_X1 U11 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  XOR2_X1 U13 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  XOR2_X1 U15 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  XOR2_X1 U17 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  XOR2_X1 U19 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  XOR2_X1 U21 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X1 U25 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  XOR2_X1 U27 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  XOR2_X1 U29 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  XOR2_X1 U31 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  XOR2_X1 U33 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  XOR2_X1 U35 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  XOR2_X1 U37 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  XOR2_X1 U39 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  XOR2_X1 U41 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  XOR2_X1 U43 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  XOR2_X1 U45 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  XOR2_X1 U47 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  XOR2_X1 U49 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  XOR2_X1 U51 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  XOR2_X1 U53 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U55 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  XOR2_X1 U57 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  XNOR2_X1 U1 ( .A(A[31]), .B(n1), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n1) );
  AND2_X1 U4 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  AND2_X1 U6 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  AND2_X1 U8 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  AND2_X1 U10 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  AND2_X1 U12 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  AND2_X1 U14 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  AND2_X1 U16 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  AND2_X1 U18 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  AND2_X1 U20 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  AND2_X1 U22 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  AND2_X1 U24 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  AND2_X1 U26 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  AND2_X1 U28 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  AND2_X1 U30 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  AND2_X1 U32 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  AND2_X1 U34 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  AND2_X1 U36 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  AND2_X1 U38 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U40 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U42 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  AND2_X1 U44 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  AND2_X1 U46 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  AND2_X1 U48 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  AND2_X1 U50 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  AND2_X1 U52 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  AND2_X1 U54 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  AND2_X1 U56 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  INV_X1 U58 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module MUX61_generic_NB32 ( A, B, C, D, E, F, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [2:0] SEL;
  output [31:0] Y;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N44, n95, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116;

  DLH_X1 \Y_reg[31]  ( .G(n115), .D(N44), .Q(Y[31]) );
  DLH_X1 \Y_reg[30]  ( .G(n115), .D(N42), .Q(Y[30]) );
  DLH_X1 \Y_reg[29]  ( .G(n114), .D(N41), .Q(Y[29]) );
  DLH_X1 \Y_reg[28]  ( .G(n115), .D(N40), .Q(Y[28]) );
  DLH_X1 \Y_reg[27]  ( .G(n115), .D(N39), .Q(Y[27]) );
  DLH_X1 \Y_reg[26]  ( .G(n115), .D(N38), .Q(Y[26]) );
  DLH_X1 \Y_reg[25]  ( .G(n115), .D(N37), .Q(Y[25]) );
  DLH_X1 \Y_reg[24]  ( .G(n115), .D(N36), .Q(Y[24]) );
  DLH_X1 \Y_reg[23]  ( .G(n115), .D(N35), .Q(Y[23]) );
  DLH_X1 \Y_reg[22]  ( .G(n115), .D(N34), .Q(Y[22]) );
  DLH_X1 \Y_reg[21]  ( .G(n115), .D(N33), .Q(Y[21]) );
  DLH_X1 \Y_reg[20]  ( .G(n116), .D(N32), .Q(Y[20]) );
  DLH_X1 \Y_reg[19]  ( .G(n116), .D(N31), .Q(Y[19]) );
  DLH_X1 \Y_reg[18]  ( .G(n116), .D(N30), .Q(Y[18]) );
  DLH_X1 \Y_reg[17]  ( .G(n116), .D(N29), .Q(Y[17]) );
  DLH_X1 \Y_reg[16]  ( .G(n116), .D(N28), .Q(Y[16]) );
  DLH_X1 \Y_reg[15]  ( .G(n116), .D(N27), .Q(Y[15]) );
  DLH_X1 \Y_reg[14]  ( .G(n116), .D(N26), .Q(Y[14]) );
  DLH_X1 \Y_reg[13]  ( .G(n116), .D(N25), .Q(Y[13]) );
  DLH_X1 \Y_reg[12]  ( .G(n116), .D(N24), .Q(Y[12]) );
  DLH_X1 \Y_reg[11]  ( .G(n115), .D(N23), .Q(Y[11]) );
  DLH_X1 \Y_reg[10]  ( .G(n116), .D(N22), .Q(Y[10]) );
  DLH_X1 \Y_reg[9]  ( .G(n114), .D(N21), .Q(Y[9]) );
  DLH_X1 \Y_reg[8]  ( .G(n114), .D(N20), .Q(Y[8]) );
  DLH_X1 \Y_reg[7]  ( .G(n114), .D(N19), .Q(Y[7]) );
  DLH_X1 \Y_reg[6]  ( .G(n114), .D(N18), .Q(Y[6]) );
  DLH_X1 \Y_reg[5]  ( .G(n114), .D(N17), .Q(Y[5]) );
  DLH_X1 \Y_reg[4]  ( .G(n114), .D(N16), .Q(Y[4]) );
  DLH_X1 \Y_reg[3]  ( .G(n114), .D(N15), .Q(Y[3]) );
  DLH_X1 \Y_reg[2]  ( .G(n114), .D(N14), .Q(Y[2]) );
  DLH_X1 \Y_reg[1]  ( .G(n114), .D(N13), .Q(Y[1]) );
  DLH_X1 \Y_reg[0]  ( .G(n114), .D(N12), .Q(Y[0]) );
  AOI222_X1 U2 ( .A1(A[25]), .A2(n99), .B1(B[25]), .B2(n104), .C1(C[25]), .C2(
        n96), .ZN(n23) );
  AOI222_X1 U3 ( .A1(A[29]), .A2(n99), .B1(B[29]), .B2(n104), .C1(C[29]), .C2(
        n96), .ZN(n15) );
  BUF_X1 U4 ( .A(n95), .Z(n114) );
  BUF_X1 U5 ( .A(n95), .Z(n115) );
  BUF_X1 U6 ( .A(n95), .Z(n116) );
  OR4_X1 U7 ( .A1(n113), .A2(n110), .A3(n107), .A4(n7), .ZN(n95) );
  OR3_X1 U8 ( .A1(n104), .A2(n99), .A3(n96), .ZN(n7) );
  BUF_X1 U9 ( .A(n5), .Z(n108) );
  BUF_X1 U10 ( .A(n5), .Z(n109) );
  BUF_X1 U11 ( .A(n9), .Z(n100) );
  BUF_X1 U12 ( .A(n10), .Z(n98) );
  BUF_X1 U13 ( .A(n6), .Z(n105) );
  BUF_X1 U14 ( .A(n8), .Z(n102) );
  BUF_X1 U15 ( .A(n6), .Z(n106) );
  BUF_X1 U16 ( .A(n4), .Z(n111) );
  BUF_X1 U17 ( .A(n4), .Z(n112) );
  BUF_X1 U18 ( .A(n6), .Z(n107) );
  BUF_X1 U19 ( .A(n9), .Z(n101) );
  BUF_X1 U20 ( .A(n4), .Z(n113) );
  BUF_X1 U21 ( .A(n9), .Z(n99) );
  BUF_X1 U22 ( .A(n5), .Z(n110) );
  BUF_X1 U23 ( .A(n10), .Z(n97) );
  BUF_X1 U24 ( .A(n8), .Z(n103) );
  BUF_X1 U25 ( .A(n10), .Z(n96) );
  BUF_X1 U26 ( .A(n8), .Z(n104) );
  NOR3_X1 U27 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n77), .ZN(n10) );
  NOR3_X1 U28 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n75), .ZN(n8) );
  NOR3_X1 U29 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n76), .ZN(n6) );
  NOR3_X1 U30 ( .A1(n75), .A2(SEL[1]), .A3(n76), .ZN(n4) );
  NOR3_X1 U31 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n9) );
  NOR3_X1 U32 ( .A1(n77), .A2(SEL[2]), .A3(n75), .ZN(n5) );
  INV_X1 U33 ( .A(SEL[0]), .ZN(n75) );
  NAND2_X1 U34 ( .A1(n49), .A2(n50), .ZN(N24) );
  AOI222_X1 U35 ( .A1(D[12]), .A2(n109), .B1(E[12]), .B2(n106), .C1(F[12]), 
        .C2(n112), .ZN(n50) );
  INV_X1 U36 ( .A(SEL[2]), .ZN(n76) );
  INV_X1 U37 ( .A(SEL[1]), .ZN(n77) );
  NAND2_X1 U38 ( .A1(n19), .A2(n20), .ZN(N39) );
  AOI222_X1 U39 ( .A1(A[27]), .A2(n99), .B1(B[27]), .B2(n104), .C1(C[27]), 
        .C2(n96), .ZN(n19) );
  AOI222_X1 U40 ( .A1(D[27]), .A2(n110), .B1(E[27]), .B2(n107), .C1(F[27]), 
        .C2(n113), .ZN(n20) );
  NAND2_X1 U41 ( .A1(n73), .A2(n74), .ZN(N12) );
  AOI222_X1 U42 ( .A1(A[0]), .A2(n101), .B1(B[0]), .B2(n102), .C1(C[0]), .C2(
        n98), .ZN(n73) );
  AOI222_X1 U43 ( .A1(D[0]), .A2(n108), .B1(E[0]), .B2(n105), .C1(F[0]), .C2(
        n111), .ZN(n74) );
  NAND2_X1 U44 ( .A1(n71), .A2(n72), .ZN(N13) );
  AOI222_X1 U45 ( .A1(A[1]), .A2(n101), .B1(B[1]), .B2(n102), .C1(C[1]), .C2(
        n98), .ZN(n71) );
  AOI222_X1 U46 ( .A1(D[1]), .A2(n108), .B1(E[1]), .B2(n105), .C1(F[1]), .C2(
        n111), .ZN(n72) );
  NAND2_X1 U47 ( .A1(n69), .A2(n70), .ZN(N14) );
  AOI222_X1 U48 ( .A1(A[2]), .A2(n101), .B1(B[2]), .B2(n102), .C1(C[2]), .C2(
        n98), .ZN(n69) );
  AOI222_X1 U49 ( .A1(D[2]), .A2(n108), .B1(E[2]), .B2(n105), .C1(F[2]), .C2(
        n111), .ZN(n70) );
  NAND2_X1 U50 ( .A1(n67), .A2(n68), .ZN(N15) );
  AOI222_X1 U51 ( .A1(A[3]), .A2(n101), .B1(B[3]), .B2(n102), .C1(C[3]), .C2(
        n98), .ZN(n67) );
  AOI222_X1 U52 ( .A1(D[3]), .A2(n108), .B1(E[3]), .B2(n105), .C1(F[3]), .C2(
        n111), .ZN(n68) );
  NAND2_X1 U53 ( .A1(n65), .A2(n66), .ZN(N16) );
  AOI222_X1 U54 ( .A1(A[4]), .A2(n101), .B1(B[4]), .B2(n102), .C1(C[4]), .C2(
        n98), .ZN(n65) );
  AOI222_X1 U55 ( .A1(D[4]), .A2(n108), .B1(E[4]), .B2(n105), .C1(F[4]), .C2(
        n111), .ZN(n66) );
  NAND2_X1 U56 ( .A1(n63), .A2(n64), .ZN(N17) );
  AOI222_X1 U57 ( .A1(A[5]), .A2(n101), .B1(B[5]), .B2(n102), .C1(C[5]), .C2(
        n98), .ZN(n63) );
  AOI222_X1 U58 ( .A1(D[5]), .A2(n108), .B1(E[5]), .B2(n105), .C1(F[5]), .C2(
        n111), .ZN(n64) );
  NAND2_X1 U59 ( .A1(n61), .A2(n62), .ZN(N18) );
  AOI222_X1 U60 ( .A1(A[6]), .A2(n101), .B1(B[6]), .B2(n102), .C1(C[6]), .C2(
        n98), .ZN(n61) );
  AOI222_X1 U61 ( .A1(D[6]), .A2(n108), .B1(E[6]), .B2(n105), .C1(F[6]), .C2(
        n111), .ZN(n62) );
  NAND2_X1 U62 ( .A1(n59), .A2(n60), .ZN(N19) );
  AOI222_X1 U63 ( .A1(A[7]), .A2(n101), .B1(B[7]), .B2(n102), .C1(C[7]), .C2(
        n98), .ZN(n59) );
  AOI222_X1 U64 ( .A1(D[7]), .A2(n108), .B1(E[7]), .B2(n105), .C1(F[7]), .C2(
        n111), .ZN(n60) );
  NAND2_X1 U65 ( .A1(n57), .A2(n58), .ZN(N20) );
  AOI222_X1 U66 ( .A1(A[8]), .A2(n101), .B1(B[8]), .B2(n102), .C1(C[8]), .C2(
        n98), .ZN(n57) );
  AOI222_X1 U67 ( .A1(D[8]), .A2(n108), .B1(E[8]), .B2(n105), .C1(F[8]), .C2(
        n111), .ZN(n58) );
  NAND2_X1 U68 ( .A1(n55), .A2(n56), .ZN(N21) );
  AOI222_X1 U69 ( .A1(A[9]), .A2(n100), .B1(B[9]), .B2(n102), .C1(C[9]), .C2(
        n97), .ZN(n55) );
  AOI222_X1 U70 ( .A1(D[9]), .A2(n108), .B1(E[9]), .B2(n105), .C1(F[9]), .C2(
        n111), .ZN(n56) );
  NAND2_X1 U71 ( .A1(n53), .A2(n54), .ZN(N22) );
  AOI222_X1 U72 ( .A1(A[10]), .A2(n100), .B1(B[10]), .B2(n102), .C1(C[10]), 
        .C2(n97), .ZN(n53) );
  AOI222_X1 U73 ( .A1(D[10]), .A2(n108), .B1(E[10]), .B2(n105), .C1(F[10]), 
        .C2(n111), .ZN(n54) );
  NAND2_X1 U74 ( .A1(n51), .A2(n52), .ZN(N23) );
  AOI222_X1 U75 ( .A1(A[11]), .A2(n100), .B1(B[11]), .B2(n102), .C1(C[11]), 
        .C2(n97), .ZN(n51) );
  AOI222_X1 U76 ( .A1(D[11]), .A2(n108), .B1(E[11]), .B2(n105), .C1(F[11]), 
        .C2(n111), .ZN(n52) );
  NAND2_X1 U77 ( .A1(n45), .A2(n46), .ZN(N26) );
  AOI222_X1 U78 ( .A1(A[14]), .A2(n100), .B1(B[14]), .B2(n103), .C1(C[14]), 
        .C2(n97), .ZN(n45) );
  AOI222_X1 U79 ( .A1(D[14]), .A2(n109), .B1(E[14]), .B2(n106), .C1(F[14]), 
        .C2(n112), .ZN(n46) );
  NAND2_X1 U80 ( .A1(n43), .A2(n44), .ZN(N27) );
  AOI222_X1 U81 ( .A1(A[15]), .A2(n100), .B1(B[15]), .B2(n103), .C1(C[15]), 
        .C2(n97), .ZN(n43) );
  AOI222_X1 U82 ( .A1(D[15]), .A2(n109), .B1(E[15]), .B2(n106), .C1(F[15]), 
        .C2(n112), .ZN(n44) );
  NAND2_X1 U83 ( .A1(n41), .A2(n42), .ZN(N28) );
  AOI222_X1 U84 ( .A1(A[16]), .A2(n100), .B1(B[16]), .B2(n103), .C1(C[16]), 
        .C2(n97), .ZN(n41) );
  AOI222_X1 U85 ( .A1(D[16]), .A2(n109), .B1(E[16]), .B2(n106), .C1(F[16]), 
        .C2(n112), .ZN(n42) );
  NAND2_X1 U86 ( .A1(n39), .A2(n40), .ZN(N29) );
  AOI222_X1 U87 ( .A1(A[17]), .A2(n100), .B1(B[17]), .B2(n103), .C1(C[17]), 
        .C2(n97), .ZN(n39) );
  AOI222_X1 U88 ( .A1(D[17]), .A2(n109), .B1(E[17]), .B2(n106), .C1(F[17]), 
        .C2(n112), .ZN(n40) );
  NAND2_X1 U89 ( .A1(n37), .A2(n38), .ZN(N30) );
  AOI222_X1 U90 ( .A1(A[18]), .A2(n100), .B1(B[18]), .B2(n103), .C1(C[18]), 
        .C2(n97), .ZN(n37) );
  AOI222_X1 U91 ( .A1(D[18]), .A2(n109), .B1(E[18]), .B2(n106), .C1(F[18]), 
        .C2(n112), .ZN(n38) );
  NAND2_X1 U92 ( .A1(n35), .A2(n36), .ZN(N31) );
  AOI222_X1 U93 ( .A1(A[19]), .A2(n100), .B1(B[19]), .B2(n103), .C1(C[19]), 
        .C2(n97), .ZN(n35) );
  AOI222_X1 U94 ( .A1(D[19]), .A2(n109), .B1(E[19]), .B2(n106), .C1(F[19]), 
        .C2(n112), .ZN(n36) );
  NAND2_X1 U95 ( .A1(n29), .A2(n30), .ZN(N34) );
  AOI222_X1 U96 ( .A1(A[22]), .A2(n99), .B1(B[22]), .B2(n103), .C1(C[22]), 
        .C2(n96), .ZN(n29) );
  AOI222_X1 U97 ( .A1(D[22]), .A2(n109), .B1(E[22]), .B2(n106), .C1(F[22]), 
        .C2(n112), .ZN(n30) );
  NAND2_X1 U98 ( .A1(n27), .A2(n28), .ZN(N35) );
  AOI222_X1 U99 ( .A1(A[23]), .A2(n99), .B1(B[23]), .B2(n103), .C1(C[23]), 
        .C2(n96), .ZN(n27) );
  AOI222_X1 U100 ( .A1(D[23]), .A2(n109), .B1(E[23]), .B2(n106), .C1(F[23]), 
        .C2(n112), .ZN(n28) );
  NAND2_X1 U101 ( .A1(n25), .A2(n26), .ZN(N36) );
  AOI222_X1 U102 ( .A1(A[24]), .A2(n99), .B1(B[24]), .B2(n104), .C1(C[24]), 
        .C2(n96), .ZN(n25) );
  AOI222_X1 U103 ( .A1(D[24]), .A2(n110), .B1(E[24]), .B2(n107), .C1(F[24]), 
        .C2(n113), .ZN(n26) );
  NAND2_X1 U104 ( .A1(n23), .A2(n24), .ZN(N37) );
  AOI222_X1 U105 ( .A1(D[25]), .A2(n110), .B1(E[25]), .B2(n107), .C1(F[25]), 
        .C2(n113), .ZN(n24) );
  NAND2_X1 U106 ( .A1(n21), .A2(n22), .ZN(N38) );
  AOI222_X1 U107 ( .A1(A[26]), .A2(n99), .B1(B[26]), .B2(n104), .C1(C[26]), 
        .C2(n96), .ZN(n21) );
  AOI222_X1 U108 ( .A1(D[26]), .A2(n110), .B1(E[26]), .B2(n107), .C1(F[26]), 
        .C2(n113), .ZN(n22) );
  NAND2_X1 U109 ( .A1(n17), .A2(n18), .ZN(N40) );
  AOI222_X1 U110 ( .A1(A[28]), .A2(n99), .B1(B[28]), .B2(n104), .C1(C[28]), 
        .C2(n96), .ZN(n17) );
  AOI222_X1 U111 ( .A1(D[28]), .A2(n110), .B1(E[28]), .B2(n107), .C1(F[28]), 
        .C2(n113), .ZN(n18) );
  NAND2_X1 U112 ( .A1(n15), .A2(n16), .ZN(N41) );
  AOI222_X1 U113 ( .A1(D[29]), .A2(n110), .B1(E[29]), .B2(n107), .C1(F[29]), 
        .C2(n113), .ZN(n16) );
  NAND2_X1 U114 ( .A1(n13), .A2(n14), .ZN(N42) );
  AOI222_X1 U115 ( .A1(A[30]), .A2(n99), .B1(B[30]), .B2(n104), .C1(C[30]), 
        .C2(n96), .ZN(n13) );
  AOI222_X1 U116 ( .A1(D[30]), .A2(n110), .B1(E[30]), .B2(n107), .C1(F[30]), 
        .C2(n113), .ZN(n14) );
  NAND2_X1 U117 ( .A1(n11), .A2(n12), .ZN(N44) );
  AOI222_X1 U118 ( .A1(A[31]), .A2(n99), .B1(B[31]), .B2(n104), .C1(C[31]), 
        .C2(n96), .ZN(n11) );
  AOI222_X1 U119 ( .A1(D[31]), .A2(n110), .B1(E[31]), .B2(n107), .C1(F[31]), 
        .C2(n113), .ZN(n12) );
  NAND2_X1 U120 ( .A1(n47), .A2(n48), .ZN(N25) );
  AOI222_X1 U121 ( .A1(A[13]), .A2(n100), .B1(B[13]), .B2(n103), .C1(C[13]), 
        .C2(n97), .ZN(n47) );
  AOI222_X1 U122 ( .A1(D[13]), .A2(n109), .B1(E[13]), .B2(n106), .C1(F[13]), 
        .C2(n112), .ZN(n48) );
  NAND2_X1 U123 ( .A1(n33), .A2(n34), .ZN(N32) );
  AOI222_X1 U124 ( .A1(A[20]), .A2(n100), .B1(B[20]), .B2(n103), .C1(C[20]), 
        .C2(n97), .ZN(n33) );
  AOI222_X1 U125 ( .A1(D[20]), .A2(n109), .B1(E[20]), .B2(n106), .C1(F[20]), 
        .C2(n112), .ZN(n34) );
  NAND2_X1 U126 ( .A1(n31), .A2(n32), .ZN(N33) );
  AOI222_X1 U127 ( .A1(A[21]), .A2(n99), .B1(B[21]), .B2(n103), .C1(C[21]), 
        .C2(n96), .ZN(n31) );
  AOI222_X1 U128 ( .A1(D[21]), .A2(n109), .B1(E[21]), .B2(n106), .C1(F[21]), 
        .C2(n112), .ZN(n32) );
  AOI222_X1 U129 ( .A1(A[12]), .A2(n100), .B1(B[12]), .B2(n103), .C1(C[12]), 
        .C2(n97), .ZN(n49) );
endmodule


module FD_NB5_0 ( CK, RESET, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module LOGIC_NB32 ( SEL, A, B, RES );
  input [3:0] SEL;
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  wire   n65, n66, n67, n69, n70, n71, n73, n74, n75, n77, n78, n79, n81, n83,
         n85, n86, n87, n89, n91, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n169,
         n170, n171, n173, n174, n175, n177, n178, n179, n181, n182, n183,
         n185, n186, n187, n189, n191, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n72, n76, n80, n82;

  AOI22_X1 U1 ( .A1(n60), .A2(n46), .B1(A[6]), .B2(n72), .ZN(n79) );
  AOI22_X1 U2 ( .A1(n63), .A2(n46), .B1(A[6]), .B2(n82), .ZN(n77) );
  AOI22_X1 U3 ( .A1(n58), .A2(n39), .B1(A[14]), .B2(n64), .ZN(n171) );
  AOI22_X1 U4 ( .A1(n61), .A2(n39), .B1(A[14]), .B2(n76), .ZN(n169) );
  AOI22_X1 U5 ( .A1(n60), .A2(n44), .B1(n72), .B2(A[9]), .ZN(n67) );
  AOI22_X1 U6 ( .A1(n63), .A2(n44), .B1(n82), .B2(A[9]), .ZN(n65) );
  BUF_X1 U7 ( .A(SEL[0]), .Z(n59) );
  BUF_X1 U8 ( .A(SEL[0]), .Z(n58) );
  OAI22_X1 U9 ( .A1(n177), .A2(n178), .B1(B[12]), .B2(n179), .ZN(RES[12]) );
  INV_X1 U10 ( .A(B[12]), .ZN(n178) );
  AOI22_X1 U11 ( .A1(n61), .A2(n41), .B1(A[12]), .B2(n76), .ZN(n177) );
  AOI22_X1 U12 ( .A1(n58), .A2(n41), .B1(A[12]), .B2(n64), .ZN(n179) );
  OAI22_X1 U13 ( .A1(n85), .A2(n86), .B1(B[4]), .B2(n87), .ZN(RES[4]) );
  INV_X1 U14 ( .A(B[4]), .ZN(n86) );
  AOI22_X1 U15 ( .A1(n63), .A2(n48), .B1(A[4]), .B2(n82), .ZN(n85) );
  AOI22_X1 U16 ( .A1(n60), .A2(n48), .B1(A[4]), .B2(n72), .ZN(n87) );
  OAI22_X1 U17 ( .A1(n101), .A2(n102), .B1(B[2]), .B2(n103), .ZN(RES[2]) );
  INV_X1 U18 ( .A(B[2]), .ZN(n102) );
  OAI22_X1 U19 ( .A1(n145), .A2(n146), .B1(B[1]), .B2(n147), .ZN(RES[1]) );
  INV_X1 U20 ( .A(B[1]), .ZN(n146) );
  AOI22_X1 U21 ( .A1(n61), .A2(n51), .B1(A[1]), .B2(n76), .ZN(n145) );
  AOI22_X1 U22 ( .A1(n58), .A2(n51), .B1(A[1]), .B2(n64), .ZN(n147) );
  OAI22_X1 U23 ( .A1(n81), .A2(n57), .B1(B[5]), .B2(n83), .ZN(RES[5]) );
  OAI22_X1 U24 ( .A1(n89), .A2(n56), .B1(B[3]), .B2(n91), .ZN(RES[3]) );
  AOI22_X1 U25 ( .A1(n63), .A2(n49), .B1(A[3]), .B2(n82), .ZN(n89) );
  AOI22_X1 U26 ( .A1(n60), .A2(n49), .B1(A[3]), .B2(n72), .ZN(n91) );
  OAI22_X1 U27 ( .A1(n73), .A2(n74), .B1(B[7]), .B2(n75), .ZN(RES[7]) );
  INV_X1 U28 ( .A(B[7]), .ZN(n74) );
  AOI22_X1 U29 ( .A1(n63), .A2(n45), .B1(A[7]), .B2(n82), .ZN(n73) );
  AOI22_X1 U30 ( .A1(n60), .A2(n45), .B1(A[7]), .B2(n72), .ZN(n75) );
  OAI22_X1 U31 ( .A1(n69), .A2(n70), .B1(B[8]), .B2(n71), .ZN(RES[8]) );
  INV_X1 U32 ( .A(B[8]), .ZN(n70) );
  AOI22_X1 U33 ( .A1(n63), .A2(n53), .B1(A[8]), .B2(n82), .ZN(n69) );
  AOI22_X1 U34 ( .A1(n60), .A2(n53), .B1(A[8]), .B2(n72), .ZN(n71) );
  OAI22_X1 U35 ( .A1(n181), .A2(n182), .B1(B[11]), .B2(n183), .ZN(RES[11]) );
  INV_X1 U36 ( .A(B[11]), .ZN(n182) );
  AOI22_X1 U37 ( .A1(n61), .A2(n42), .B1(A[11]), .B2(n76), .ZN(n181) );
  AOI22_X1 U38 ( .A1(n58), .A2(n42), .B1(A[11]), .B2(n64), .ZN(n183) );
  OAI22_X1 U39 ( .A1(n173), .A2(n174), .B1(B[13]), .B2(n175), .ZN(RES[13]) );
  INV_X1 U40 ( .A(B[13]), .ZN(n174) );
  OAI22_X1 U41 ( .A1(n165), .A2(n166), .B1(B[15]), .B2(n167), .ZN(RES[15]) );
  INV_X1 U42 ( .A(B[15]), .ZN(n166) );
  AOI22_X1 U43 ( .A1(n61), .A2(n52), .B1(A[15]), .B2(n76), .ZN(n165) );
  AOI22_X1 U44 ( .A1(n58), .A2(n52), .B1(A[15]), .B2(n64), .ZN(n167) );
  OAI22_X1 U45 ( .A1(n93), .A2(n94), .B1(B[31]), .B2(n95), .ZN(RES[31]) );
  INV_X1 U46 ( .A(B[31]), .ZN(n94) );
  AOI22_X1 U47 ( .A1(n63), .A2(n96), .B1(A[31]), .B2(n82), .ZN(n93) );
  AOI22_X1 U48 ( .A1(n60), .A2(n96), .B1(A[31]), .B2(n72), .ZN(n95) );
  OAI22_X1 U49 ( .A1(n185), .A2(n186), .B1(B[10]), .B2(n187), .ZN(RES[10]) );
  INV_X1 U50 ( .A(B[10]), .ZN(n186) );
  AOI22_X1 U51 ( .A1(n61), .A2(n43), .B1(A[10]), .B2(n76), .ZN(n185) );
  AOI22_X1 U52 ( .A1(n58), .A2(n43), .B1(A[10]), .B2(n64), .ZN(n187) );
  OAI22_X1 U53 ( .A1(n157), .A2(n158), .B1(B[17]), .B2(n159), .ZN(RES[17]) );
  INV_X1 U54 ( .A(B[17]), .ZN(n158) );
  AOI22_X1 U55 ( .A1(n61), .A2(n160), .B1(A[17]), .B2(n76), .ZN(n157) );
  AOI22_X1 U56 ( .A1(n58), .A2(n160), .B1(A[17]), .B2(n64), .ZN(n159) );
  OAI22_X1 U57 ( .A1(n153), .A2(n154), .B1(B[18]), .B2(n155), .ZN(RES[18]) );
  INV_X1 U58 ( .A(B[18]), .ZN(n154) );
  AOI22_X1 U59 ( .A1(n61), .A2(n156), .B1(A[18]), .B2(n76), .ZN(n153) );
  AOI22_X1 U60 ( .A1(n58), .A2(n156), .B1(A[18]), .B2(n64), .ZN(n155) );
  OAI22_X1 U61 ( .A1(n161), .A2(n162), .B1(B[16]), .B2(n163), .ZN(RES[16]) );
  INV_X1 U62 ( .A(B[16]), .ZN(n162) );
  AOI22_X1 U63 ( .A1(n61), .A2(n164), .B1(A[16]), .B2(n76), .ZN(n161) );
  AOI22_X1 U64 ( .A1(n58), .A2(n164), .B1(A[16]), .B2(n64), .ZN(n163) );
  OAI22_X1 U65 ( .A1(n117), .A2(n118), .B1(B[26]), .B2(n119), .ZN(RES[26]) );
  INV_X1 U66 ( .A(B[26]), .ZN(n118) );
  AOI22_X1 U67 ( .A1(n62), .A2(n120), .B1(A[26]), .B2(n80), .ZN(n117) );
  AOI22_X1 U68 ( .A1(n59), .A2(n120), .B1(A[26]), .B2(n68), .ZN(n119) );
  OAI22_X1 U69 ( .A1(n133), .A2(n134), .B1(B[22]), .B2(n135), .ZN(RES[22]) );
  INV_X1 U70 ( .A(B[22]), .ZN(n134) );
  AOI22_X1 U71 ( .A1(n62), .A2(n136), .B1(A[22]), .B2(n80), .ZN(n133) );
  AOI22_X1 U72 ( .A1(n59), .A2(n136), .B1(A[22]), .B2(n68), .ZN(n135) );
  OAI22_X1 U73 ( .A1(n97), .A2(n98), .B1(B[30]), .B2(n99), .ZN(RES[30]) );
  INV_X1 U74 ( .A(B[30]), .ZN(n98) );
  AOI22_X1 U75 ( .A1(n62), .A2(n100), .B1(A[30]), .B2(n80), .ZN(n97) );
  AOI22_X1 U76 ( .A1(n59), .A2(n100), .B1(A[30]), .B2(n68), .ZN(n99) );
  OAI22_X1 U77 ( .A1(n121), .A2(n122), .B1(B[25]), .B2(n123), .ZN(RES[25]) );
  INV_X1 U78 ( .A(B[25]), .ZN(n122) );
  AOI22_X1 U79 ( .A1(n62), .A2(n124), .B1(A[25]), .B2(n80), .ZN(n121) );
  AOI22_X1 U80 ( .A1(n59), .A2(n124), .B1(A[25]), .B2(n68), .ZN(n123) );
  OAI22_X1 U81 ( .A1(n109), .A2(n110), .B1(B[28]), .B2(n111), .ZN(RES[28]) );
  INV_X1 U82 ( .A(B[28]), .ZN(n110) );
  AOI22_X1 U83 ( .A1(n62), .A2(n112), .B1(A[28]), .B2(n80), .ZN(n109) );
  AOI22_X1 U84 ( .A1(n59), .A2(n112), .B1(A[28]), .B2(n68), .ZN(n111) );
  OAI22_X1 U85 ( .A1(n137), .A2(n138), .B1(B[21]), .B2(n139), .ZN(RES[21]) );
  INV_X1 U86 ( .A(B[21]), .ZN(n138) );
  AOI22_X1 U87 ( .A1(n62), .A2(n140), .B1(A[21]), .B2(n80), .ZN(n137) );
  AOI22_X1 U88 ( .A1(n59), .A2(n140), .B1(A[21]), .B2(n68), .ZN(n139) );
  OAI22_X1 U89 ( .A1(n125), .A2(n126), .B1(B[24]), .B2(n127), .ZN(RES[24]) );
  INV_X1 U90 ( .A(B[24]), .ZN(n126) );
  AOI22_X1 U91 ( .A1(n62), .A2(n128), .B1(A[24]), .B2(n80), .ZN(n125) );
  AOI22_X1 U92 ( .A1(n59), .A2(n128), .B1(A[24]), .B2(n68), .ZN(n127) );
  OAI22_X1 U93 ( .A1(n113), .A2(n114), .B1(B[27]), .B2(n115), .ZN(RES[27]) );
  INV_X1 U94 ( .A(B[27]), .ZN(n114) );
  AOI22_X1 U95 ( .A1(n62), .A2(n116), .B1(A[27]), .B2(n80), .ZN(n113) );
  AOI22_X1 U96 ( .A1(n59), .A2(n116), .B1(A[27]), .B2(n68), .ZN(n115) );
  OAI22_X1 U97 ( .A1(n129), .A2(n130), .B1(B[23]), .B2(n131), .ZN(RES[23]) );
  INV_X1 U98 ( .A(B[23]), .ZN(n130) );
  AOI22_X1 U99 ( .A1(n62), .A2(n132), .B1(A[23]), .B2(n80), .ZN(n129) );
  AOI22_X1 U100 ( .A1(n59), .A2(n132), .B1(A[23]), .B2(n68), .ZN(n131) );
  OAI22_X1 U101 ( .A1(n105), .A2(n106), .B1(B[29]), .B2(n107), .ZN(RES[29]) );
  INV_X1 U102 ( .A(B[29]), .ZN(n106) );
  AOI22_X1 U103 ( .A1(n62), .A2(n108), .B1(A[29]), .B2(n80), .ZN(n105) );
  AOI22_X1 U104 ( .A1(n59), .A2(n108), .B1(A[29]), .B2(n68), .ZN(n107) );
  OAI22_X1 U105 ( .A1(n141), .A2(n142), .B1(B[20]), .B2(n143), .ZN(RES[20]) );
  INV_X1 U106 ( .A(B[20]), .ZN(n142) );
  AOI22_X1 U107 ( .A1(n62), .A2(n144), .B1(A[20]), .B2(n80), .ZN(n141) );
  AOI22_X1 U108 ( .A1(n59), .A2(n144), .B1(A[20]), .B2(n68), .ZN(n143) );
  OAI22_X1 U109 ( .A1(n149), .A2(n150), .B1(B[19]), .B2(n151), .ZN(RES[19]) );
  INV_X1 U110 ( .A(B[19]), .ZN(n150) );
  AOI22_X1 U111 ( .A1(n61), .A2(n152), .B1(A[19]), .B2(n76), .ZN(n149) );
  AOI22_X1 U112 ( .A1(n58), .A2(n152), .B1(A[19]), .B2(n64), .ZN(n151) );
  BUF_X1 U113 ( .A(SEL[0]), .Z(n60) );
  INV_X1 U114 ( .A(A[31]), .ZN(n96) );
  INV_X1 U115 ( .A(A[17]), .ZN(n160) );
  INV_X1 U116 ( .A(A[18]), .ZN(n156) );
  INV_X1 U117 ( .A(A[16]), .ZN(n164) );
  INV_X1 U118 ( .A(A[26]), .ZN(n120) );
  INV_X1 U119 ( .A(A[22]), .ZN(n136) );
  INV_X1 U120 ( .A(A[30]), .ZN(n100) );
  INV_X1 U121 ( .A(A[27]), .ZN(n116) );
  INV_X1 U122 ( .A(A[23]), .ZN(n132) );
  INV_X1 U123 ( .A(A[29]), .ZN(n108) );
  INV_X1 U124 ( .A(A[19]), .ZN(n152) );
  INV_X1 U125 ( .A(A[25]), .ZN(n124) );
  INV_X1 U126 ( .A(A[28]), .ZN(n112) );
  INV_X1 U127 ( .A(A[21]), .ZN(n140) );
  INV_X1 U128 ( .A(A[24]), .ZN(n128) );
  INV_X1 U129 ( .A(A[20]), .ZN(n144) );
  BUF_X1 U130 ( .A(SEL[1]), .Z(n62) );
  BUF_X1 U131 ( .A(SEL[1]), .Z(n61) );
  BUF_X1 U132 ( .A(SEL[2]), .Z(n68) );
  BUF_X1 U133 ( .A(SEL[3]), .Z(n80) );
  BUF_X1 U134 ( .A(SEL[2]), .Z(n64) );
  BUF_X1 U135 ( .A(SEL[3]), .Z(n76) );
  BUF_X1 U136 ( .A(SEL[2]), .Z(n72) );
  BUF_X1 U137 ( .A(SEL[3]), .Z(n82) );
  BUF_X1 U138 ( .A(SEL[1]), .Z(n63) );
  INV_X1 U139 ( .A(A[14]), .ZN(n39) );
  INV_X1 U140 ( .A(A[13]), .ZN(n40) );
  INV_X1 U141 ( .A(A[12]), .ZN(n41) );
  INV_X1 U142 ( .A(A[11]), .ZN(n42) );
  INV_X1 U143 ( .A(A[10]), .ZN(n43) );
  INV_X1 U144 ( .A(A[9]), .ZN(n44) );
  INV_X1 U145 ( .A(A[7]), .ZN(n45) );
  INV_X1 U146 ( .A(A[6]), .ZN(n46) );
  INV_X1 U147 ( .A(A[5]), .ZN(n47) );
  INV_X1 U148 ( .A(A[4]), .ZN(n48) );
  INV_X1 U149 ( .A(A[3]), .ZN(n49) );
  INV_X1 U150 ( .A(A[2]), .ZN(n50) );
  INV_X1 U151 ( .A(A[1]), .ZN(n51) );
  OAI22_X1 U152 ( .A1(n189), .A2(n55), .B1(B[0]), .B2(n191), .ZN(RES[0]) );
  OAI22_X1 U153 ( .A1(n77), .A2(n78), .B1(B[6]), .B2(n79), .ZN(RES[6]) );
  INV_X1 U154 ( .A(B[6]), .ZN(n78) );
  OAI22_X1 U155 ( .A1(n169), .A2(n170), .B1(B[14]), .B2(n171), .ZN(RES[14]) );
  INV_X1 U156 ( .A(B[14]), .ZN(n170) );
  AOI22_X1 U157 ( .A1(n61), .A2(n40), .B1(A[13]), .B2(n76), .ZN(n173) );
  AOI22_X1 U158 ( .A1(n58), .A2(n40), .B1(A[13]), .B2(n64), .ZN(n175) );
  AOI22_X1 U159 ( .A1(n59), .A2(n50), .B1(A[2]), .B2(n68), .ZN(n103) );
  AOI22_X1 U160 ( .A1(n62), .A2(n50), .B1(A[2]), .B2(n80), .ZN(n101) );
  AOI22_X1 U161 ( .A1(n63), .A2(n47), .B1(A[5]), .B2(n82), .ZN(n81) );
  AOI22_X1 U162 ( .A1(n60), .A2(n47), .B1(A[5]), .B2(n72), .ZN(n83) );
  OAI22_X1 U163 ( .A1(n65), .A2(n66), .B1(B[9]), .B2(n67), .ZN(RES[9]) );
  INV_X1 U164 ( .A(B[9]), .ZN(n66) );
  AOI22_X1 U165 ( .A1(n61), .A2(n54), .B1(A[0]), .B2(n76), .ZN(n189) );
  AOI22_X1 U166 ( .A1(n58), .A2(n54), .B1(A[0]), .B2(n64), .ZN(n191) );
  INV_X1 U167 ( .A(A[15]), .ZN(n52) );
  INV_X1 U168 ( .A(A[8]), .ZN(n53) );
  INV_X1 U169 ( .A(A[0]), .ZN(n54) );
  INV_X1 U170 ( .A(B[0]), .ZN(n55) );
  INV_X1 U171 ( .A(B[3]), .ZN(n56) );
  INV_X1 U172 ( .A(B[5]), .ZN(n57) );
endmodule


module COMPARATOR_NB32 ( AdderRes, MSB, CO, OP_CODE, US, SOUT );
  input [31:0] AdderRes;
  input [1:0] MSB;
  input [2:0] OP_CODE;
  output [31:0] SOUT;
  input CO, US;
  wire   n6, n7, n8, n9, n10, n13, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n3, n4, n5;
  assign SOUT[31] = 1'b0;
  assign SOUT[30] = 1'b0;
  assign SOUT[29] = 1'b0;
  assign SOUT[28] = 1'b0;
  assign SOUT[27] = 1'b0;
  assign SOUT[26] = 1'b0;
  assign SOUT[25] = 1'b0;
  assign SOUT[24] = 1'b0;
  assign SOUT[23] = 1'b0;
  assign SOUT[22] = 1'b0;
  assign SOUT[21] = 1'b0;
  assign SOUT[20] = 1'b0;
  assign SOUT[19] = 1'b0;
  assign SOUT[18] = 1'b0;
  assign SOUT[17] = 1'b0;
  assign SOUT[16] = 1'b0;
  assign SOUT[15] = 1'b0;
  assign SOUT[14] = 1'b0;
  assign SOUT[13] = 1'b0;
  assign SOUT[12] = 1'b0;
  assign SOUT[11] = 1'b0;
  assign SOUT[10] = 1'b0;
  assign SOUT[9] = 1'b0;
  assign SOUT[8] = 1'b0;
  assign SOUT[7] = 1'b0;
  assign SOUT[6] = 1'b0;
  assign SOUT[5] = 1'b0;
  assign SOUT[4] = 1'b0;
  assign SOUT[3] = 1'b0;
  assign SOUT[2] = 1'b0;
  assign SOUT[1] = 1'b0;

  NAND3_X1 U29 ( .A1(n4), .A2(n5), .A3(n13), .ZN(n10) );
  INV_X1 U2 ( .A(n15), .ZN(n19) );
  NOR4_X1 U3 ( .A1(AdderRes[1]), .A2(AdderRes[19]), .A3(AdderRes[18]), .A4(
        AdderRes[17]), .ZN(n27) );
  NOR2_X1 U4 ( .A1(n23), .A2(n24), .ZN(n15) );
  NAND4_X1 U5 ( .A1(n29), .A2(n30), .A3(n31), .A4(n32), .ZN(n23) );
  NAND4_X1 U6 ( .A1(n25), .A2(n26), .A3(n27), .A4(n28), .ZN(n24) );
  NOR4_X1 U7 ( .A1(AdderRes[9]), .A2(AdderRes[8]), .A3(AdderRes[7]), .A4(
        AdderRes[6]), .ZN(n32) );
  AOI211_X1 U8 ( .C1(OP_CODE[0]), .C2(n15), .A(n5), .B(n4), .ZN(n17) );
  OAI221_X1 U9 ( .B1(n6), .B2(n7), .C1(n8), .C2(n9), .A(n10), .ZN(SOUT[0]) );
  INV_X1 U10 ( .A(n9), .ZN(n7) );
  AOI22_X1 U11 ( .A1(n16), .A2(OP_CODE[2]), .B1(CO), .B2(n17), .ZN(n8) );
  XNOR2_X1 U12 ( .A(n3), .B(n15), .ZN(n13) );
  AND2_X1 U13 ( .A1(n4), .A2(n18), .ZN(n16) );
  OAI21_X1 U14 ( .B1(n19), .B2(OP_CODE[0]), .A(CO), .ZN(n18) );
  AOI22_X1 U15 ( .A1(n21), .A2(MSB[1]), .B1(MSB[0]), .B2(n17), .ZN(n6) );
  NOR2_X1 U16 ( .A1(OP_CODE[1]), .A2(n22), .ZN(n21) );
  AOI22_X1 U17 ( .A1(OP_CODE[0]), .A2(n19), .B1(OP_CODE[2]), .B2(n3), .ZN(n22)
         );
  NOR2_X1 U18 ( .A1(US), .A2(n20), .ZN(n9) );
  XNOR2_X1 U19 ( .A(MSB[0]), .B(MSB[1]), .ZN(n20) );
  INV_X1 U20 ( .A(OP_CODE[0]), .ZN(n3) );
  NOR4_X1 U21 ( .A1(AdderRes[12]), .A2(AdderRes[11]), .A3(AdderRes[10]), .A4(
        AdderRes[0]), .ZN(n25) );
  NOR4_X1 U22 ( .A1(AdderRes[5]), .A2(AdderRes[4]), .A3(AdderRes[3]), .A4(
        AdderRes[31]), .ZN(n31) );
  NOR4_X1 U23 ( .A1(AdderRes[27]), .A2(AdderRes[26]), .A3(AdderRes[25]), .A4(
        AdderRes[24]), .ZN(n29) );
  NOR4_X1 U24 ( .A1(AdderRes[16]), .A2(AdderRes[15]), .A3(AdderRes[14]), .A4(
        AdderRes[13]), .ZN(n26) );
  NOR4_X1 U25 ( .A1(AdderRes[30]), .A2(AdderRes[2]), .A3(AdderRes[29]), .A4(
        AdderRes[28]), .ZN(n30) );
  NOR4_X1 U26 ( .A1(AdderRes[23]), .A2(AdderRes[22]), .A3(AdderRes[21]), .A4(
        AdderRes[20]), .ZN(n28) );
  INV_X1 U27 ( .A(OP_CODE[1]), .ZN(n4) );
  INV_X1 U28 ( .A(OP_CODE[2]), .ZN(n5) );
endmodule


module SHIFTER_NB32_LS5 ( FUNC, US, DATA1, DATA2, OUTSHFT );
  input [1:0] FUNC;
  input [31:0] DATA1;
  input [4:0] DATA2;
  output [31:0] OUTSHFT;
  input US;
  wire   n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n349, n350, n351, n353, n355, n356, n357, n358, n359, n360,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n586, n588, n590, n591, n592, n593, n594, n595, n596,
         n599, n600, n601, n603, n604, n605, n608, n609, n611, n614, n615,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n628, n630,
         n632, n633, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n172, n290, n348, n352, n354, n361, n557, n585, n587, n589,
         n597, n598, n602, n606, n607, n610, n612, n613, n616, n617, n627,
         n629, n631, n634, n657, n669, n680, n719, n735, n736, n737, n738,
         n739;

  NAND3_X1 U608 ( .A1(n221), .A2(n738), .A3(n151), .ZN(n220) );
  NAND3_X1 U609 ( .A1(n255), .A2(n256), .A3(n257), .ZN(OUTSHFT[30]) );
  NAND3_X1 U610 ( .A1(n282), .A2(n283), .A3(n284), .ZN(OUTSHFT[29]) );
  NAND3_X1 U611 ( .A1(n303), .A2(n162), .A3(n138), .ZN(n302) );
  NAND3_X1 U612 ( .A1(n309), .A2(n310), .A3(n311), .ZN(OUTSHFT[27]) );
  NAND3_X1 U613 ( .A1(n322), .A2(n323), .A3(n324), .ZN(OUTSHFT[26]) );
  NAND3_X1 U614 ( .A1(n335), .A2(n336), .A3(n337), .ZN(OUTSHFT[25]) );
  NAND3_X1 U615 ( .A1(n398), .A2(n399), .A3(n400), .ZN(OUTSHFT[23]) );
  NAND3_X1 U616 ( .A1(n422), .A2(n423), .A3(n424), .ZN(OUTSHFT[22]) );
  NAND3_X1 U617 ( .A1(n221), .A2(n738), .A3(n260), .ZN(n472) );
  NAND3_X1 U618 ( .A1(n502), .A2(n503), .A3(n504), .ZN(OUTSHFT[19]) );
  NAND3_X1 U619 ( .A1(n520), .A2(n521), .A3(n522), .ZN(OUTSHFT[18]) );
  NAND3_X1 U620 ( .A1(n532), .A2(n533), .A3(n534), .ZN(OUTSHFT[17]) );
  NAND3_X1 U621 ( .A1(DATA2[4]), .A2(FUNC[0]), .A3(FUNC[1]), .ZN(n552) );
  NAND3_X1 U622 ( .A1(FUNC[0]), .A2(n254), .A3(FUNC[1]), .ZN(n301) );
  AOI221_X1 U2 ( .B1(n121), .B2(DATA1[17]), .C1(n118), .C2(DATA1[18]), .A(n726), .ZN(n385) );
  AOI221_X1 U3 ( .B1(n121), .B2(DATA1[27]), .C1(DATA1[26]), .C2(n118), .A(n718), .ZN(n397) );
  AOI221_X1 U4 ( .B1(DATA1[26]), .B2(n121), .C1(n118), .C2(DATA1[27]), .A(n599), .ZN(n363) );
  AOI221_X1 U5 ( .B1(n121), .B2(DATA1[8]), .C1(n118), .C2(DATA1[7]), .A(n615), 
        .ZN(n367) );
  AOI221_X1 U6 ( .B1(n121), .B2(DATA1[17]), .C1(n118), .C2(DATA1[16]), .A(n705), .ZN(n440) );
  AOI221_X1 U7 ( .B1(n111), .B2(DATA1[26]), .C1(DATA1[25]), .C2(n103), .A(n695), .ZN(n445) );
  AOI221_X1 U8 ( .B1(n121), .B2(DATA1[24]), .C1(DATA1[25]), .C2(n118), .A(n663), .ZN(n405) );
  NAND2_X1 U9 ( .A1(n251), .A2(n254), .ZN(n148) );
  AND2_X1 U10 ( .A1(n738), .A2(n641), .ZN(n87) );
  AOI221_X1 U11 ( .B1(n121), .B2(DATA1[3]), .C1(n118), .C2(DATA1[2]), .A(n724), 
        .ZN(n394) );
  AOI221_X1 U12 ( .B1(n121), .B2(DATA1[6]), .C1(n118), .C2(DATA1[5]), .A(n670), 
        .ZN(n414) );
  INV_X1 U13 ( .A(n361), .ZN(n142) );
  INV_X1 U14 ( .A(n135), .ZN(n128) );
  INV_X1 U15 ( .A(n361), .ZN(n143) );
  INV_X1 U16 ( .A(n136), .ZN(n129) );
  INV_X1 U17 ( .A(n126), .ZN(n124) );
  INV_X1 U18 ( .A(n126), .ZN(n125) );
  INV_X1 U19 ( .A(n108), .ZN(n104) );
  INV_X1 U20 ( .A(n108), .ZN(n103) );
  INV_X1 U21 ( .A(n617), .ZN(n589) );
  OAI21_X1 U22 ( .B1(n413), .B2(n358), .A(n512), .ZN(n238) );
  INV_X1 U23 ( .A(n617), .ZN(n597) );
  INV_X1 U24 ( .A(n278), .ZN(n272) );
  BUF_X1 U25 ( .A(n87), .Z(n134) );
  BUF_X1 U26 ( .A(n87), .Z(n135) );
  BUF_X1 U27 ( .A(n141), .Z(n361) );
  BUF_X1 U28 ( .A(n138), .Z(n136) );
  BUF_X1 U29 ( .A(n87), .Z(n137) );
  INV_X1 U30 ( .A(n427), .ZN(n219) );
  BUF_X1 U31 ( .A(n138), .Z(n130) );
  BUF_X1 U32 ( .A(n138), .Z(n131) );
  BUF_X1 U33 ( .A(n87), .Z(n132) );
  BUF_X1 U34 ( .A(n87), .Z(n133) );
  BUF_X1 U35 ( .A(n139), .Z(n144) );
  BUF_X1 U36 ( .A(n139), .Z(n145) );
  BUF_X1 U37 ( .A(n139), .Z(n146) );
  BUF_X1 U38 ( .A(n140), .Z(n290) );
  BUF_X1 U39 ( .A(n140), .Z(n172) );
  BUF_X1 U40 ( .A(n140), .Z(n348) );
  BUF_X1 U41 ( .A(n141), .Z(n352) );
  BUF_X1 U42 ( .A(n141), .Z(n354) );
  INV_X1 U43 ( .A(n344), .ZN(n456) );
  NAND2_X1 U44 ( .A1(n512), .A2(n219), .ZN(n228) );
  INV_X1 U45 ( .A(n212), .ZN(n463) );
  INV_X1 U46 ( .A(n325), .ZN(n687) );
  BUF_X1 U47 ( .A(n87), .Z(n138) );
  NOR3_X1 U48 ( .A1(n698), .A2(n711), .A3(n699), .ZN(n278) );
  OAI222_X1 U49 ( .A1(n506), .A2(n361), .B1(n408), .B2(n128), .C1(n678), .C2(
        n616), .ZN(n318) );
  INV_X1 U50 ( .A(n412), .ZN(n678) );
  INV_X1 U51 ( .A(n118), .ZN(n117) );
  INV_X1 U52 ( .A(n115), .ZN(n110) );
  NOR2_X1 U53 ( .A1(n633), .A2(n609), .ZN(n344) );
  OAI221_X1 U54 ( .B1(n390), .B2(n172), .C1(n391), .C2(n124), .A(n378), .ZN(
        n178) );
  OAI21_X1 U55 ( .B1(n120), .B2(n246), .A(n278), .ZN(n447) );
  OAI22_X1 U56 ( .A1(n483), .A2(n128), .B1(n647), .B2(n598), .ZN(n640) );
  OAI22_X1 U57 ( .A1(n288), .A2(n598), .B1(n347), .B2(n128), .ZN(n159) );
  OAI22_X1 U58 ( .A1(n278), .A2(n598), .B1(n435), .B2(n129), .ZN(n198) );
  NOR2_X1 U59 ( .A1(n124), .A2(n246), .ZN(n427) );
  AOI22_X1 U60 ( .A1(n688), .A2(n589), .B1(n450), .B2(n131), .ZN(n328) );
  AOI22_X1 U61 ( .A1(n170), .A2(n265), .B1(n629), .B2(n176), .ZN(n374) );
  BUF_X1 U62 ( .A(n153), .Z(n634) );
  AOI21_X1 U63 ( .B1(n426), .B2(n142), .A(n427), .ZN(n196) );
  INV_X1 U64 ( .A(n428), .ZN(n426) );
  BUF_X1 U65 ( .A(n153), .Z(n657) );
  NOR3_X1 U66 ( .A1(n556), .A2(n112), .A3(n129), .ZN(n555) );
  OAI21_X1 U67 ( .B1(n468), .B2(n122), .A(n537), .ZN(n500) );
  OAI21_X1 U68 ( .B1(n263), .B2(n144), .A(n438), .ZN(n200) );
  OAI21_X1 U69 ( .B1(n278), .B2(n144), .A(n690), .ZN(n330) );
  OAI21_X1 U70 ( .B1(n288), .B2(n145), .A(n464), .ZN(n212) );
  OAI21_X1 U71 ( .B1(n364), .B2(n123), .A(n603), .ZN(n294) );
  OAI21_X1 U72 ( .B1(n576), .B2(n358), .A(n571), .ZN(n268) );
  INV_X1 U73 ( .A(n447), .ZN(n576) );
  OAI21_X1 U74 ( .B1(n288), .B2(n122), .A(n537), .ZN(n492) );
  OAI21_X1 U75 ( .B1(n344), .B2(n123), .A(n603), .ZN(n286) );
  OAI21_X1 U76 ( .B1(n278), .B2(n358), .A(n571), .ZN(n261) );
  OAI21_X1 U77 ( .B1(n263), .B2(n122), .A(n527), .ZN(n276) );
  OAI21_X1 U78 ( .B1(n428), .B2(n128), .A(n315), .ZN(n259) );
  INV_X1 U79 ( .A(n116), .ZN(n111) );
  OAI21_X1 U80 ( .B1(n354), .B2(n248), .A(n406), .ZN(n188) );
  OAI21_X1 U81 ( .B1(n428), .B2(n602), .A(n343), .ZN(n325) );
  OAI21_X1 U82 ( .B1(n428), .B2(n123), .A(n527), .ZN(n277) );
  OAI21_X1 U83 ( .B1(n344), .B2(n144), .A(n346), .ZN(n152) );
  NAND2_X1 U84 ( .A1(n260), .A2(n130), .ZN(n507) );
  NAND2_X1 U85 ( .A1(n289), .A2(n131), .ZN(n247) );
  BUF_X1 U86 ( .A(n109), .Z(n108) );
  INV_X1 U87 ( .A(n265), .ZN(n548) );
  BUF_X1 U88 ( .A(n587), .Z(n616) );
  INV_X1 U89 ( .A(n540), .ZN(n350) );
  INV_X1 U90 ( .A(n530), .ZN(n441) );
  BUF_X1 U91 ( .A(n557), .Z(n598) );
  BUF_X1 U92 ( .A(n109), .Z(n105) );
  BUF_X1 U93 ( .A(n109), .Z(n106) );
  INV_X1 U94 ( .A(n248), .ZN(n655) );
  INV_X1 U95 ( .A(n263), .ZN(n688) );
  BUF_X1 U96 ( .A(n109), .Z(n107) );
  BUF_X1 U97 ( .A(n557), .Z(n602) );
  INV_X1 U98 ( .A(n516), .ZN(n413) );
  INV_X1 U99 ( .A(n480), .ZN(n390) );
  BUF_X1 U100 ( .A(n585), .Z(n607) );
  BUF_X1 U101 ( .A(n557), .Z(n606) );
  BUF_X1 U102 ( .A(n585), .Z(n610) );
  BUF_X1 U103 ( .A(n585), .Z(n612) );
  BUF_X1 U104 ( .A(n587), .Z(n613) );
  INV_X1 U105 ( .A(n185), .ZN(n404) );
  INV_X1 U106 ( .A(n467), .ZN(n364) );
  BUF_X1 U107 ( .A(n587), .Z(n617) );
  INV_X1 U108 ( .A(n369), .ZN(n468) );
  INV_X1 U109 ( .A(n179), .ZN(n401) );
  INV_X1 U110 ( .A(n376), .ZN(n174) );
  INV_X1 U111 ( .A(n334), .ZN(n333) );
  INV_X1 U112 ( .A(n513), .ZN(n512) );
  OAI21_X1 U113 ( .B1(n514), .B2(n145), .A(n515), .ZN(n513) );
  INV_X1 U114 ( .A(n298), .ZN(n635) );
  INV_X1 U115 ( .A(n316), .ZN(n313) );
  INV_X1 U116 ( .A(n156), .ZN(n155) );
  AOI22_X1 U117 ( .A1(n157), .A2(n158), .B1(n159), .B2(n160), .ZN(n156) );
  INV_X1 U118 ( .A(n582), .ZN(n580) );
  AOI22_X1 U119 ( .A1(n286), .A2(n151), .B1(n291), .B2(n634), .ZN(n582) );
  INV_X1 U120 ( .A(n568), .ZN(n566) );
  AOI22_X1 U121 ( .A1(n261), .A2(n151), .B1(n264), .B2(n634), .ZN(n568) );
  INV_X1 U122 ( .A(n210), .ZN(n208) );
  BUF_X1 U123 ( .A(n345), .Z(n139) );
  BUF_X1 U124 ( .A(n345), .Z(n141) );
  BUF_X1 U125 ( .A(n345), .Z(n140) );
  INV_X1 U126 ( .A(n340), .ZN(n338) );
  AOI22_X1 U127 ( .A1(n152), .A2(n260), .B1(n157), .B2(n258), .ZN(n340) );
  AOI221_X1 U128 ( .B1(n121), .B2(DATA1[7]), .C1(n118), .C2(DATA1[6]), .A(n723), .ZN(n395) );
  OAI22_X1 U129 ( .A1(n98), .A2(n113), .B1(n97), .B2(n107), .ZN(n723) );
  NAND2_X1 U130 ( .A1(n148), .A2(n186), .ZN(n265) );
  AOI221_X1 U131 ( .B1(n121), .B2(DATA1[10]), .C1(n118), .C2(DATA1[9]), .A(
        n668), .ZN(n418) );
  OAI22_X1 U132 ( .A1(n95), .A2(n113), .B1(n680), .B2(n106), .ZN(n668) );
  AOI222_X1 U133 ( .A1(n451), .A2(n589), .B1(n443), .B2(n133), .C1(n450), .C2(
        n142), .ZN(n527) );
  AOI222_X1 U134 ( .A1(n371), .A2(n142), .B1(n353), .B2(n589), .C1(n471), .C2(
        n133), .ZN(n537) );
  OAI222_X1 U135 ( .A1(n396), .A2(n354), .B1(n397), .B2(n616), .C1(n485), .C2(
        n129), .ZN(n216) );
  INV_X1 U136 ( .A(n383), .ZN(n485) );
  AOI21_X1 U137 ( .B1(n118), .B2(n102), .A(n604), .ZN(n288) );
  OAI221_X1 U138 ( .B1(n119), .B2(n98), .C1(n117), .C2(n97), .A(n679), .ZN(
        n412) );
  AOI22_X1 U139 ( .A1(DATA1[7]), .A2(n111), .B1(DATA1[6]), .B2(n103), .ZN(n679) );
  OAI221_X1 U140 ( .B1(n119), .B2(n95), .C1(n586), .C2(n680), .A(n709), .ZN(
        n434) );
  AOI22_X1 U141 ( .A1(DATA1[10]), .A2(n110), .B1(DATA1[9]), .B2(n104), .ZN(
        n709) );
  AOI222_X1 U142 ( .A1(n366), .A2(n142), .B1(n460), .B2(n133), .C1(n365), .C2(
        n589), .ZN(n603) );
  AOI222_X1 U143 ( .A1(n449), .A2(n142), .B1(n433), .B2(n133), .C1(n434), .C2(
        n589), .ZN(n571) );
  AOI221_X1 U144 ( .B1(n387), .B2(n136), .C1(n388), .C2(n597), .A(n730), .ZN(
        n547) );
  OAI22_X1 U145 ( .A1(n146), .A2(n647), .B1(n125), .B2(n642), .ZN(n730) );
  OAI222_X1 U146 ( .A1(n395), .A2(n361), .B1(n394), .B2(n616), .C1(n379), .C2(
        n358), .ZN(n304) );
  AOI21_X1 U147 ( .B1(n590), .B2(n102), .A(n689), .ZN(n263) );
  OAI221_X1 U148 ( .B1(n584), .B2(n611), .C1(n117), .C2(n246), .A(n344), .ZN(
        n467) );
  OAI221_X1 U149 ( .B1(n120), .B2(n100), .C1(n586), .C2(n101), .A(n666), .ZN(
        n516) );
  NOR2_X1 U150 ( .A1(n633), .A2(n655), .ZN(n666) );
  AOI221_X1 U151 ( .B1(n402), .B2(n127), .C1(n403), .C2(n142), .A(n404), .ZN(
        n179) );
  INV_X1 U152 ( .A(n405), .ZN(n402) );
  AOI221_X1 U153 ( .B1(n447), .B2(n142), .C1(n448), .C2(n127), .A(n707), .ZN(
        n334) );
  INV_X1 U154 ( .A(n690), .ZN(n707) );
  OAI221_X1 U155 ( .B1(n119), .B2(n600), .C1(n586), .C2(n611), .A(n729), .ZN(
        n480) );
  AOI21_X1 U156 ( .B1(n102), .B2(n103), .A(n713), .ZN(n729) );
  AOI221_X1 U157 ( .B1(n392), .B2(n135), .C1(n478), .C2(n126), .A(n479), .ZN(
        n213) );
  OAI22_X1 U158 ( .A1(n613), .A2(n390), .B1(n146), .B2(n391), .ZN(n479) );
  AOI221_X1 U159 ( .B1(n480), .B2(n136), .C1(n650), .C2(n589), .A(n725), .ZN(
        n543) );
  OAI22_X1 U160 ( .A1(n146), .A2(n384), .B1(n125), .B2(n385), .ZN(n725) );
  INV_X1 U161 ( .A(n329), .ZN(n289) );
  OAI221_X1 U162 ( .B1(n468), .B2(n290), .C1(n469), .C2(n124), .A(n464), .ZN(
        n211) );
  INV_X1 U163 ( .A(n370), .ZN(n469) );
  OAI221_X1 U164 ( .B1(n367), .B2(n352), .C1(n350), .C2(n125), .A(n605), .ZN(
        n293) );
  AOI22_X1 U165 ( .A1(n135), .A2(n369), .B1(n597), .B2(n370), .ZN(n605) );
  AOI21_X1 U166 ( .B1(n115), .B2(n102), .A(n689), .ZN(n428) );
  OAI221_X1 U167 ( .B1(n528), .B2(n122), .C1(n441), .C2(n146), .A(n572), .ZN(
        n267) );
  AOI22_X1 U168 ( .A1(n134), .A2(n573), .B1(n597), .B2(n439), .ZN(n572) );
  OAI221_X1 U169 ( .B1(n347), .B2(n128), .C1(n367), .C2(n124), .A(n368), .ZN(
        n164) );
  AOI22_X1 U170 ( .A1(n589), .A2(n369), .B1(n142), .B2(n370), .ZN(n368) );
  OAI221_X1 U171 ( .B1(n436), .B2(n172), .C1(n437), .C2(n124), .A(n438), .ZN(
        n199) );
  INV_X1 U172 ( .A(n439), .ZN(n437) );
  OAI221_X1 U173 ( .B1(n413), .B2(n290), .C1(n414), .C2(n124), .A(n406), .ZN(
        n187) );
  OAI221_X1 U174 ( .B1(n394), .B2(n172), .C1(n395), .C2(n124), .A(n174), .ZN(
        n177) );
  OAI221_X1 U175 ( .B1(n574), .B2(n129), .C1(n441), .C2(n125), .A(n696), .ZN(
        n331) );
  AOI22_X1 U176 ( .A1(n589), .A2(n573), .B1(n143), .B2(n439), .ZN(n696) );
  OAI221_X1 U177 ( .B1(n508), .B2(n125), .C1(n405), .C2(n610), .A(n558), .ZN(
        n252) );
  AOI22_X1 U178 ( .A1(n143), .A2(n559), .B1(n137), .B2(n403), .ZN(n558) );
  OAI221_X1 U179 ( .B1(n584), .B2(n91), .C1(n117), .C2(n92), .A(n614), .ZN(
        n540) );
  AOI22_X1 U180 ( .A1(DATA1[9]), .A2(n110), .B1(DATA1[10]), .B2(n103), .ZN(
        n614) );
  OAI221_X1 U181 ( .B1(n584), .B2(n94), .C1(n117), .C2(n680), .A(n700), .ZN(
        n530) );
  AOI22_X1 U182 ( .A1(DATA1[6]), .A2(n111), .B1(DATA1[7]), .B2(n103), .ZN(n700) );
  OAI221_X1 U183 ( .B1(n483), .B2(n348), .C1(n385), .C2(n128), .A(n484), .ZN(
        n217) );
  AOI22_X1 U184 ( .A1(n126), .A2(n393), .B1(n597), .B2(n387), .ZN(n484) );
  OAI221_X1 U185 ( .B1(n363), .B2(n358), .C1(n364), .C2(n145), .A(n346), .ZN(
        n165) );
  OAI221_X1 U186 ( .B1(n445), .B2(n352), .C1(n429), .C2(n125), .A(n531), .ZN(
        n281) );
  AOI22_X1 U187 ( .A1(n134), .A2(n447), .B1(n597), .B2(n448), .ZN(n531) );
  OAI221_X1 U188 ( .B1(n445), .B2(n123), .C1(n435), .C2(n128), .A(n446), .ZN(
        n201) );
  AOI22_X1 U189 ( .A1(n589), .A2(n447), .B1(n142), .B2(n448), .ZN(n446) );
  OAI221_X1 U190 ( .B1(n405), .B2(n348), .C1(n407), .C2(n124), .A(n519), .ZN(
        n239) );
  AOI22_X1 U191 ( .A1(n134), .A2(n235), .B1(n597), .B2(n403), .ZN(n519) );
  OAI221_X1 U192 ( .B1(n457), .B2(n123), .C1(n363), .C2(n610), .A(n541), .ZN(
        n501) );
  AOI22_X1 U193 ( .A1(n143), .A2(n542), .B1(n138), .B2(n467), .ZN(n541) );
  OAI221_X1 U194 ( .B1(n405), .B2(n128), .C1(n407), .C2(n612), .A(n656), .ZN(
        n320) );
  AOI22_X1 U195 ( .A1(n143), .A2(n410), .B1(n127), .B2(n411), .ZN(n656) );
  OAI221_X1 U196 ( .B1(n395), .B2(n129), .C1(n379), .C2(n606), .A(n481), .ZN(
        n222) );
  AOI22_X1 U197 ( .A1(n142), .A2(n482), .B1(n127), .B2(n382), .ZN(n481) );
  OAI221_X1 U198 ( .B1(n384), .B2(n128), .C1(n385), .C2(n602), .A(n386), .ZN(
        n170) );
  AOI22_X1 U199 ( .A1(n142), .A2(n387), .B1(n127), .B2(n388), .ZN(n386) );
  OAI221_X1 U200 ( .B1(n356), .B2(n129), .C1(n357), .C2(n125), .A(n359), .ZN(
        n154) );
  AOI22_X1 U201 ( .A1(n589), .A2(n360), .B1(n143), .B2(n362), .ZN(n359) );
  OAI221_X1 U202 ( .B1(n440), .B2(n290), .C1(n441), .C2(n128), .A(n442), .ZN(
        n193) );
  AOI22_X1 U203 ( .A1(n127), .A2(n443), .B1(n597), .B2(n444), .ZN(n442) );
  INV_X1 U204 ( .A(n455), .ZN(n260) );
  OAI221_X1 U205 ( .B1(n528), .B2(n128), .C1(n440), .C2(n613), .A(n702), .ZN(
        n332) );
  AOI22_X1 U206 ( .A1(n143), .A2(n443), .B1(n126), .B2(n451), .ZN(n702) );
  OAI221_X1 U207 ( .B1(n414), .B2(n129), .C1(n418), .C2(n607), .A(n517), .ZN(
        n233) );
  AOI22_X1 U208 ( .A1(n143), .A2(n421), .B1(n126), .B2(n518), .ZN(n517) );
  OAI221_X1 U209 ( .B1(n538), .B2(n358), .C1(n367), .C2(n607), .A(n539), .ZN(
        n489) );
  AOI22_X1 U210 ( .A1(n143), .A2(n540), .B1(n137), .B2(n370), .ZN(n539) );
  OAI221_X1 U211 ( .B1(n458), .B2(n129), .C1(n357), .C2(n607), .A(n536), .ZN(
        n499) );
  AOI22_X1 U212 ( .A1(n126), .A2(n366), .B1(n142), .B2(n365), .ZN(n536) );
  OAI221_X1 U213 ( .B1(n524), .B2(n129), .C1(n525), .C2(n607), .A(n526), .ZN(
        n279) );
  INV_X1 U214 ( .A(n433), .ZN(n525) );
  AOI22_X1 U215 ( .A1(n126), .A2(n449), .B1(n143), .B2(n434), .ZN(n526) );
  OAI221_X1 U216 ( .B1(n508), .B2(n129), .C1(n509), .C2(n606), .A(n510), .ZN(
        n237) );
  AOI22_X1 U217 ( .A1(n142), .A2(n511), .B1(n127), .B2(n412), .ZN(n510) );
  OAI221_X1 U218 ( .B1(n528), .B2(n352), .C1(n440), .C2(n124), .A(n529), .ZN(
        n273) );
  AOI22_X1 U219 ( .A1(n589), .A2(n530), .B1(n136), .B2(n439), .ZN(n529) );
  OAI221_X1 U220 ( .B1(n417), .B2(n348), .C1(n418), .C2(n128), .A(n419), .ZN(
        n183) );
  AOI22_X1 U221 ( .A1(n126), .A2(n420), .B1(n597), .B2(n421), .ZN(n419) );
  OAI221_X1 U222 ( .B1(n440), .B2(n129), .C1(n574), .C2(n125), .A(n575), .ZN(
        n266) );
  AOI22_X1 U223 ( .A1(n589), .A2(n443), .B1(n142), .B2(n451), .ZN(n575) );
  OAI221_X1 U224 ( .B1(n394), .B2(n129), .C1(n395), .C2(n613), .A(n720), .ZN(
        n550) );
  AOI22_X1 U225 ( .A1(n142), .A2(n643), .B1(n127), .B2(n482), .ZN(n720) );
  OAI221_X1 U226 ( .B1(n379), .B2(n128), .C1(n380), .C2(n606), .A(n381), .ZN(
        n176) );
  AOI22_X1 U227 ( .A1(n142), .A2(n382), .B1(n126), .B2(n383), .ZN(n381) );
  OAI221_X1 U228 ( .B1(n671), .B2(n129), .C1(n417), .C2(n610), .A(n672), .ZN(
        n321) );
  INV_X1 U229 ( .A(n421), .ZN(n671) );
  AOI22_X1 U230 ( .A1(n143), .A2(n420), .B1(n126), .B2(n416), .ZN(n672) );
  OAI221_X1 U231 ( .B1(n538), .B2(n129), .C1(n349), .C2(n612), .A(n618), .ZN(
        n292) );
  AOI22_X1 U232 ( .A1(n143), .A2(n353), .B1(n126), .B2(n371), .ZN(n618) );
  OAI221_X1 U233 ( .B1(n349), .B2(n172), .C1(n350), .C2(n129), .A(n351), .ZN(
        n161) );
  AOI22_X1 U234 ( .A1(n126), .A2(n353), .B1(n597), .B2(n355), .ZN(n351) );
  OAI221_X1 U235 ( .B1(n414), .B2(n348), .C1(n418), .C2(n125), .A(n665), .ZN(
        n312) );
  AOI22_X1 U236 ( .A1(n135), .A2(n415), .B1(n597), .B2(n516), .ZN(n665) );
  OAI221_X1 U237 ( .B1(n509), .B2(n129), .C1(n408), .C2(n610), .A(n561), .ZN(
        n253) );
  AOI22_X1 U238 ( .A1(n127), .A2(n235), .B1(n143), .B2(n412), .ZN(n561) );
  OAI221_X1 U239 ( .B1(n397), .B2(n354), .C1(n396), .C2(n125), .A(n714), .ZN(
        n549) );
  AOI22_X1 U240 ( .A1(n135), .A2(n382), .B1(n597), .B2(n383), .ZN(n714) );
  OAI221_X1 U241 ( .B1(n385), .B2(n352), .C1(n391), .C2(n128), .A(n649), .ZN(
        n298) );
  AOI22_X1 U242 ( .A1(n127), .A2(n387), .B1(n597), .B2(n478), .ZN(n649) );
  OAI221_X1 U243 ( .B1(n414), .B2(n616), .C1(n418), .C2(n145), .A(n562), .ZN(
        n242) );
  AOI22_X1 U244 ( .A1(n126), .A2(n421), .B1(n137), .B2(n516), .ZN(n562) );
  OAI221_X1 U245 ( .B1(n367), .B2(n128), .C1(n350), .C2(n606), .A(n470), .ZN(
        n206) );
  AOI22_X1 U246 ( .A1(n142), .A2(n355), .B1(n127), .B2(n471), .ZN(n470) );
  OAI221_X1 U247 ( .B1(n445), .B2(n129), .C1(n429), .C2(n613), .A(n691), .ZN(
        n326) );
  AOI22_X1 U248 ( .A1(n143), .A2(n432), .B1(n127), .B2(n433), .ZN(n691) );
  OAI221_X1 U249 ( .B1(n457), .B2(n128), .C1(n458), .C2(n602), .A(n459), .ZN(
        n205) );
  AOI22_X1 U250 ( .A1(n142), .A2(n460), .B1(n127), .B2(n365), .ZN(n459) );
  OAI221_X1 U251 ( .B1(n429), .B2(n128), .C1(n430), .C2(n124), .A(n431), .ZN(
        n192) );
  INV_X1 U252 ( .A(n434), .ZN(n430) );
  AOI22_X1 U253 ( .A1(n589), .A2(n432), .B1(n143), .B2(n433), .ZN(n431) );
  OAI221_X1 U254 ( .B1(n380), .B2(n128), .C1(n397), .C2(n125), .A(n648), .ZN(
        n306) );
  AOI22_X1 U255 ( .A1(n143), .A2(n383), .B1(n597), .B2(n382), .ZN(n648) );
  OAI221_X1 U256 ( .B1(n417), .B2(n129), .C1(n514), .C2(n125), .A(n560), .ZN(
        n241) );
  AOI22_X1 U257 ( .A1(n589), .A2(n420), .B1(n143), .B2(n416), .ZN(n560) );
  OAI221_X1 U258 ( .B1(n363), .B2(n129), .C1(n356), .C2(n612), .A(n583), .ZN(
        n291) );
  AOI22_X1 U259 ( .A1(n143), .A2(n360), .B1(n127), .B2(n362), .ZN(n583) );
  OAI221_X1 U260 ( .B1(n524), .B2(n122), .C1(n445), .C2(n612), .A(n569), .ZN(
        n264) );
  AOI22_X1 U261 ( .A1(n143), .A2(n570), .B1(n137), .B2(n448), .ZN(n569) );
  OAI221_X1 U262 ( .B1(n407), .B2(n128), .C1(n408), .C2(n124), .A(n409), .ZN(
        n182) );
  AOI22_X1 U263 ( .A1(n589), .A2(n410), .B1(n142), .B2(n411), .ZN(n409) );
  AOI221_X1 U264 ( .B1(n638), .B2(n136), .C1(n627), .C2(n304), .A(n639), .ZN(
        n637) );
  AND2_X1 U265 ( .A1(n303), .A2(n644), .ZN(n638) );
  OAI22_X1 U266 ( .A1(n305), .A2(n186), .B1(n197), .B2(n315), .ZN(n639) );
  NOR2_X1 U267 ( .A1(n186), .A2(n129), .ZN(n236) );
  INV_X1 U268 ( .A(n314), .ZN(n258) );
  OAI22_X1 U269 ( .A1(n396), .A2(n598), .B1(n397), .B2(n128), .ZN(n376) );
  OAI22_X1 U270 ( .A1(n108), .A2(n611), .B1(n115), .B2(n600), .ZN(n604) );
  OAI21_X1 U271 ( .B1(n119), .B2(n719), .A(n288), .ZN(n369) );
  OAI221_X1 U272 ( .B1(n547), .B2(n462), .C1(n543), .C2(n148), .A(n712), .ZN(
        OUTSHFT[0]) );
  AOI222_X1 U273 ( .A1(n550), .A2(n162), .B1(n236), .B2(n713), .C1(n644), .C2(
        n549), .ZN(n712) );
  AOI22_X1 U274 ( .A1(n371), .A2(n597), .B1(n353), .B2(n132), .ZN(n464) );
  AOI22_X1 U275 ( .A1(n450), .A2(n589), .B1(n451), .B2(n132), .ZN(n438) );
  AOI22_X1 U276 ( .A1(n415), .A2(n589), .B1(n416), .B2(n131), .ZN(n406) );
  AOI22_X1 U277 ( .A1(n392), .A2(n597), .B1(n393), .B2(n131), .ZN(n378) );
  AOI22_X1 U278 ( .A1(n365), .A2(n130), .B1(n366), .B2(n589), .ZN(n346) );
  NOR2_X1 U279 ( .A1(n245), .A2(n254), .ZN(n227) );
  AOI22_X1 U280 ( .A1(n434), .A2(n130), .B1(n449), .B2(n597), .ZN(n690) );
  AOI22_X1 U281 ( .A1(n412), .A2(n130), .B1(n235), .B2(n589), .ZN(n185) );
  AOI22_X1 U282 ( .A1(n416), .A2(n597), .B1(n420), .B2(n132), .ZN(n515) );
  AOI22_X1 U283 ( .A1(n456), .A2(n597), .B1(n366), .B2(n132), .ZN(n209) );
  INV_X1 U284 ( .A(n175), .ZN(n160) );
  NOR2_X1 U285 ( .A1(n611), .A2(n115), .ZN(n689) );
  INV_X1 U286 ( .A(n186), .ZN(n151) );
  OAI22_X1 U287 ( .A1(n738), .A2(n173), .B1(n174), .B2(n175), .ZN(n171) );
  OAI22_X1 U288 ( .A1(n195), .A2(n186), .B1(n196), .B2(n197), .ZN(n194) );
  INV_X1 U289 ( .A(n198), .ZN(n195) );
  AOI21_X1 U290 ( .B1(n221), .B2(n737), .A(n640), .ZN(n305) );
  AOI21_X1 U291 ( .B1(n403), .B2(n127), .A(n318), .ZN(n316) );
  NOR3_X1 U292 ( .A1(n175), .A2(n288), .A3(n128), .ZN(n581) );
  NOR3_X1 U293 ( .A1(n175), .A2(n263), .A3(n129), .ZN(n567) );
  AOI22_X1 U294 ( .A1(n306), .A2(n162), .B1(n645), .B2(n307), .ZN(n636) );
  INV_X1 U295 ( .A(n148), .ZN(n645) );
  BUF_X1 U296 ( .A(n163), .Z(n629) );
  OAI21_X1 U297 ( .B1(n314), .B2(n315), .A(n173), .ZN(n308) );
  OAI21_X1 U298 ( .B1(n738), .B2(n319), .A(n515), .ZN(n230) );
  OAI21_X1 U299 ( .B1(n436), .B2(n122), .A(n527), .ZN(n280) );
  OAI21_X1 U300 ( .B1(n314), .B2(n343), .A(n173), .ZN(n389) );
  OAI21_X1 U301 ( .B1(n394), .B2(n123), .A(n477), .ZN(n223) );
  INV_X1 U302 ( .A(n216), .ZN(n477) );
  OAI21_X1 U303 ( .B1(n354), .B2(n377), .A(n378), .ZN(n169) );
  OAI21_X1 U304 ( .B1(n341), .B2(n129), .A(n315), .ZN(n285) );
  BUF_X1 U305 ( .A(n163), .Z(n627) );
  OAI21_X1 U306 ( .B1(n341), .B2(n144), .A(n219), .ZN(n210) );
  NAND2_X1 U307 ( .A1(n102), .A2(n128), .ZN(n315) );
  OAI21_X1 U308 ( .B1(n341), .B2(n602), .A(n343), .ZN(n157) );
  OAI21_X1 U309 ( .B1(n341), .B2(n123), .A(n537), .ZN(n493) );
  OAI211_X1 U310 ( .C1(n486), .C2(n148), .A(n487), .B(n488), .ZN(OUTSHFT[1])
         );
  INV_X1 U311 ( .A(n501), .ZN(n486) );
  AOI22_X1 U312 ( .A1(n634), .A2(n499), .B1(n629), .B2(n500), .ZN(n487) );
  AOI221_X1 U313 ( .B1(n236), .B2(n456), .C1(n489), .C2(n234), .A(n490), .ZN(
        n488) );
  OAI211_X1 U314 ( .C1(n269), .C2(n148), .A(n270), .B(n271), .ZN(OUTSHFT[2])
         );
  INV_X1 U315 ( .A(n281), .ZN(n269) );
  AOI22_X1 U316 ( .A1(n634), .A2(n279), .B1(n631), .B2(n280), .ZN(n270) );
  AOI221_X1 U317 ( .B1(n236), .B2(n272), .C1(n273), .C2(n234), .A(n274), .ZN(
        n271) );
  OAI211_X1 U318 ( .C1(n224), .C2(n148), .A(n225), .B(n226), .ZN(OUTSHFT[3])
         );
  INV_X1 U319 ( .A(n239), .ZN(n224) );
  AOI22_X1 U320 ( .A1(n634), .A2(n237), .B1(n631), .B2(n238), .ZN(n225) );
  AOI221_X1 U321 ( .B1(n227), .B2(n228), .C1(n229), .C2(n230), .A(n231), .ZN(
        n226) );
  OAI211_X1 U322 ( .C1(n213), .C2(n148), .A(n214), .B(n215), .ZN(OUTSHFT[4])
         );
  AOI22_X1 U323 ( .A1(n222), .A2(n162), .B1(n631), .B2(n223), .ZN(n214) );
  AOI221_X1 U324 ( .B1(n160), .B2(n216), .C1(n634), .C2(n217), .A(n218), .ZN(
        n215) );
  OAI21_X1 U325 ( .B1(n197), .B2(n219), .A(n220), .ZN(n218) );
  OAI211_X1 U326 ( .C1(n202), .C2(n148), .A(n203), .B(n204), .ZN(OUTSHFT[5])
         );
  AOI22_X1 U327 ( .A1(n627), .A2(n211), .B1(n160), .B2(n212), .ZN(n203) );
  AOI221_X1 U328 ( .B1(n634), .B2(n205), .C1(n206), .C2(n162), .A(n207), .ZN(
        n204) );
  OAI22_X1 U329 ( .A1(n208), .A2(n197), .B1(n209), .B2(n186), .ZN(n207) );
  OAI211_X1 U330 ( .C1(n189), .C2(n148), .A(n190), .B(n191), .ZN(OUTSHFT[6])
         );
  INV_X1 U331 ( .A(n201), .ZN(n189) );
  AOI22_X1 U332 ( .A1(n627), .A2(n199), .B1(n160), .B2(n200), .ZN(n190) );
  AOI221_X1 U333 ( .B1(n634), .B2(n192), .C1(n193), .C2(n162), .A(n194), .ZN(
        n191) );
  OAI211_X1 U334 ( .C1(n179), .C2(n148), .A(n180), .B(n181), .ZN(OUTSHFT[7])
         );
  AOI22_X1 U335 ( .A1(n627), .A2(n187), .B1(n160), .B2(n188), .ZN(n180) );
  AOI221_X1 U336 ( .B1(n634), .B2(n182), .C1(n183), .C2(n162), .A(n184), .ZN(
        n181) );
  OAI22_X1 U337 ( .A1(n738), .A2(n173), .B1(n185), .B2(n186), .ZN(n184) );
  OAI211_X1 U338 ( .C1(n166), .C2(n148), .A(n167), .B(n168), .ZN(OUTSHFT[8])
         );
  INV_X1 U339 ( .A(n178), .ZN(n166) );
  AOI22_X1 U340 ( .A1(n176), .A2(n162), .B1(n631), .B2(n177), .ZN(n167) );
  AOI221_X1 U341 ( .B1(n151), .B2(n169), .C1(n657), .C2(n170), .A(n171), .ZN(
        n168) );
  OAI211_X1 U342 ( .C1(n147), .C2(n148), .A(n149), .B(n150), .ZN(OUTSHFT[9])
         );
  INV_X1 U343 ( .A(n165), .ZN(n147) );
  AOI22_X1 U344 ( .A1(n161), .A2(n162), .B1(n629), .B2(n164), .ZN(n149) );
  AOI221_X1 U345 ( .B1(n151), .B2(n152), .C1(n657), .C2(n154), .A(n155), .ZN(
        n150) );
  OAI211_X1 U346 ( .C1(n334), .C2(n148), .A(n684), .B(n685), .ZN(OUTSHFT[10])
         );
  AOI22_X1 U347 ( .A1(n332), .A2(n162), .B1(n629), .B2(n331), .ZN(n684) );
  AOI221_X1 U348 ( .B1(n634), .B2(n326), .C1(n151), .C2(n330), .A(n686), .ZN(
        n685) );
  OAI22_X1 U349 ( .A1(n687), .A2(n197), .B1(n328), .B2(n175), .ZN(n686) );
  OAI211_X1 U350 ( .C1(n316), .C2(n148), .A(n651), .B(n652), .ZN(OUTSHFT[11])
         );
  AOI22_X1 U351 ( .A1(n321), .A2(n162), .B1(n629), .B2(n312), .ZN(n651) );
  AOI221_X1 U352 ( .B1(n151), .B2(n318), .C1(n657), .C2(n320), .A(n653), .ZN(
        n652) );
  OAI21_X1 U353 ( .B1(n197), .B2(n315), .A(n654), .ZN(n653) );
  OAI211_X1 U354 ( .C1(n577), .C2(n148), .A(n578), .B(n579), .ZN(OUTSHFT[13])
         );
  INV_X1 U355 ( .A(n294), .ZN(n577) );
  AOI22_X1 U356 ( .A1(n292), .A2(n162), .B1(n629), .B2(n293), .ZN(n578) );
  AOI211_X1 U357 ( .C1(n158), .C2(n285), .A(n580), .B(n581), .ZN(n579) );
  OAI211_X1 U358 ( .C1(n563), .C2(n148), .A(n564), .B(n565), .ZN(OUTSHFT[14])
         );
  INV_X1 U359 ( .A(n268), .ZN(n563) );
  AOI22_X1 U360 ( .A1(n266), .A2(n162), .B1(n629), .B2(n267), .ZN(n564) );
  AOI211_X1 U361 ( .C1(n158), .C2(n259), .A(n566), .B(n567), .ZN(n565) );
  NOR2_X1 U362 ( .A1(n100), .A2(n115), .ZN(n698) );
  NOR2_X1 U363 ( .A1(n719), .A2(n586), .ZN(n699) );
  NOR2_X1 U364 ( .A1(n719), .A2(n105), .ZN(n633) );
  OAI21_X1 U365 ( .B1(n278), .B2(n507), .A(n173), .ZN(n523) );
  INV_X1 U366 ( .A(n102), .ZN(n246) );
  NAND4_X1 U367 ( .A1(n472), .A2(n173), .A3(n473), .A4(n474), .ZN(OUTSHFT[20])
         );
  AOI22_X1 U368 ( .A1(n258), .A2(n427), .B1(n289), .B2(n216), .ZN(n473) );
  AOI221_X1 U369 ( .B1(n217), .B2(n265), .C1(n629), .C2(n222), .A(n475), .ZN(
        n474) );
  OAI211_X1 U370 ( .C1(n543), .C2(n462), .A(n544), .B(n545), .ZN(OUTSHFT[16])
         );
  INV_X1 U371 ( .A(n546), .ZN(n545) );
  AOI22_X1 U372 ( .A1(n549), .A2(n162), .B1(n629), .B2(n550), .ZN(n544) );
  OAI221_X1 U373 ( .B1(n547), .B2(n548), .C1(n507), .C2(n377), .A(n173), .ZN(
        n546) );
  NOR2_X1 U374 ( .A1(n101), .A2(n105), .ZN(n711) );
  NOR2_X1 U375 ( .A1(n101), .A2(n114), .ZN(n609) );
  NAND2_X1 U376 ( .A1(n737), .A2(n102), .ZN(n343) );
  OAI21_X1 U377 ( .B1(n209), .B2(n455), .A(n173), .ZN(n454) );
  OAI21_X1 U378 ( .B1(n288), .B2(n247), .A(n173), .ZN(n287) );
  OAI21_X1 U379 ( .B1(n196), .B2(n314), .A(n173), .ZN(n425) );
  OAI21_X1 U380 ( .B1(n344), .B2(n507), .A(n173), .ZN(n535) );
  OAI21_X1 U381 ( .B1(n506), .B2(n507), .A(n173), .ZN(n505) );
  OAI21_X1 U382 ( .B1(n263), .B2(n247), .A(n173), .ZN(n262) );
  OAI21_X1 U383 ( .B1(n328), .B2(n329), .A(n173), .ZN(n327) );
  INV_X1 U384 ( .A(n574), .ZN(n450) );
  NAND2_X1 U385 ( .A1(n102), .A2(n110), .ZN(n248) );
  NAND4_X1 U386 ( .A1(n372), .A2(n373), .A3(n374), .A4(n375), .ZN(OUTSHFT[24])
         );
  INV_X1 U387 ( .A(n389), .ZN(n373) );
  AOI22_X1 U388 ( .A1(n243), .A2(n177), .B1(n657), .B2(n178), .ZN(n372) );
  AOI22_X1 U389 ( .A1(n289), .A2(n376), .B1(n260), .B2(n169), .ZN(n375) );
  INV_X1 U390 ( .A(n444), .ZN(n528) );
  INV_X1 U391 ( .A(n197), .ZN(n158) );
  INV_X1 U392 ( .A(n235), .ZN(n506) );
  BUF_X1 U393 ( .A(n88), .Z(n115) );
  INV_X1 U394 ( .A(n518), .ZN(n417) );
  INV_X1 U395 ( .A(n650), .ZN(n391) );
  NOR2_X1 U396 ( .A1(n737), .A2(n319), .ZN(n317) );
  INV_X1 U397 ( .A(n643), .ZN(n379) );
  NAND2_X1 U398 ( .A1(n737), .A2(n641), .ZN(n345) );
  INV_X1 U399 ( .A(n377), .ZN(n713) );
  INV_X1 U400 ( .A(n586), .ZN(n118) );
  AOI22_X1 U401 ( .A1(n317), .A2(n289), .B1(n260), .B2(n318), .ZN(n310) );
  AOI22_X1 U402 ( .A1(n320), .A2(n265), .B1(n629), .B2(n321), .ZN(n309) );
  AOI221_X1 U403 ( .B1(n243), .B2(n312), .C1(n634), .C2(n313), .A(n308), .ZN(
        n311) );
  INV_X1 U404 ( .A(n542), .ZN(n356) );
  INV_X1 U405 ( .A(n570), .ZN(n429) );
  INV_X1 U406 ( .A(n559), .ZN(n407) );
  INV_X1 U407 ( .A(n511), .ZN(n408) );
  INV_X1 U408 ( .A(n436), .ZN(n573) );
  BUF_X1 U409 ( .A(n163), .Z(n631) );
  INV_X1 U410 ( .A(n303), .ZN(n396) );
  BUF_X1 U411 ( .A(n88), .Z(n116) );
  INV_X1 U412 ( .A(n371), .ZN(n347) );
  INV_X1 U413 ( .A(n392), .ZN(n642) );
  AOI22_X1 U414 ( .A1(n627), .A2(n183), .B1(n243), .B2(n187), .ZN(n398) );
  AOI22_X1 U415 ( .A1(n260), .A2(n404), .B1(n182), .B2(n265), .ZN(n399) );
  AOI221_X1 U416 ( .B1(n289), .B2(n188), .C1(n657), .C2(n401), .A(n389), .ZN(
        n400) );
  AOI22_X1 U417 ( .A1(n289), .A2(n492), .B1(n657), .B2(n501), .ZN(n532) );
  AOI22_X1 U418 ( .A1(n627), .A2(n489), .B1(n243), .B2(n500), .ZN(n533) );
  AOI221_X1 U419 ( .B1(n258), .B2(n493), .C1(n499), .C2(n265), .A(n535), .ZN(
        n534) );
  AOI22_X1 U420 ( .A1(n289), .A2(n276), .B1(n657), .B2(n281), .ZN(n520) );
  AOI22_X1 U421 ( .A1(n627), .A2(n273), .B1(n243), .B2(n280), .ZN(n521) );
  AOI221_X1 U422 ( .B1(n258), .B2(n277), .C1(n279), .C2(n265), .A(n523), .ZN(
        n522) );
  AOI22_X1 U423 ( .A1(n289), .A2(n230), .B1(n657), .B2(n239), .ZN(n502) );
  AOI22_X1 U424 ( .A1(n627), .A2(n233), .B1(n243), .B2(n238), .ZN(n503) );
  AOI221_X1 U425 ( .B1(n258), .B2(n228), .C1(n237), .C2(n265), .A(n505), .ZN(
        n504) );
  AOI22_X1 U426 ( .A1(n289), .A2(n200), .B1(n657), .B2(n201), .ZN(n422) );
  AOI22_X1 U427 ( .A1(n627), .A2(n193), .B1(n243), .B2(n199), .ZN(n423) );
  AOI221_X1 U428 ( .B1(n260), .B2(n198), .C1(n192), .C2(n265), .A(n425), .ZN(
        n424) );
  AOI22_X1 U429 ( .A1(n260), .A2(n330), .B1(n243), .B2(n331), .ZN(n323) );
  AOI22_X1 U430 ( .A1(n627), .A2(n332), .B1(n657), .B2(n333), .ZN(n322) );
  AOI221_X1 U431 ( .B1(n258), .B2(n325), .C1(n326), .C2(n265), .A(n327), .ZN(
        n324) );
  INV_X1 U432 ( .A(n415), .ZN(n514) );
  AOI22_X1 U433 ( .A1(n243), .A2(n293), .B1(n657), .B2(n294), .ZN(n282) );
  AOI22_X1 U434 ( .A1(n291), .A2(n265), .B1(n629), .B2(n292), .ZN(n283) );
  AOI221_X1 U435 ( .B1(n258), .B2(n285), .C1(n260), .C2(n286), .A(n287), .ZN(
        n284) );
  AOI22_X1 U436 ( .A1(n243), .A2(n267), .B1(n657), .B2(n268), .ZN(n255) );
  AOI22_X1 U437 ( .A1(n264), .A2(n265), .B1(n631), .B2(n266), .ZN(n256) );
  AOI221_X1 U438 ( .B1(n258), .B2(n259), .C1(n260), .C2(n261), .A(n262), .ZN(
        n257) );
  INV_X1 U439 ( .A(n449), .ZN(n435) );
  BUF_X1 U440 ( .A(n88), .Z(n112) );
  BUF_X1 U441 ( .A(n88), .Z(n113) );
  BUF_X1 U442 ( .A(n358), .Z(n123) );
  BUF_X1 U443 ( .A(n358), .Z(n122) );
  BUF_X1 U444 ( .A(n88), .Z(n114) );
  INV_X1 U445 ( .A(n410), .ZN(n508) );
  INV_X1 U446 ( .A(n360), .ZN(n457) );
  INV_X1 U447 ( .A(n432), .ZN(n524) );
  INV_X1 U448 ( .A(n355), .ZN(n538) );
  INV_X1 U449 ( .A(n478), .ZN(n384) );
  INV_X1 U450 ( .A(n482), .ZN(n380) );
  INV_X1 U451 ( .A(n411), .ZN(n509) );
  INV_X1 U452 ( .A(n362), .ZN(n458) );
  INV_X1 U453 ( .A(n388), .ZN(n483) );
  INV_X1 U454 ( .A(n393), .ZN(n647) );
  INV_X1 U455 ( .A(n471), .ZN(n349) );
  INV_X1 U456 ( .A(n460), .ZN(n357) );
  NAND2_X1 U457 ( .A1(n160), .A2(n102), .ZN(n556) );
  INV_X1 U458 ( .A(n462), .ZN(n153) );
  INV_X1 U459 ( .A(n646), .ZN(n307) );
  AOI221_X1 U460 ( .B1(n392), .B2(n143), .C1(n480), .C2(n127), .A(n640), .ZN(
        n646) );
  NAND2_X1 U461 ( .A1(n295), .A2(n296), .ZN(OUTSHFT[28]) );
  AOI221_X1 U462 ( .B1(n627), .B2(n306), .C1(n634), .C2(n307), .A(n308), .ZN(
        n295) );
  AOI221_X1 U463 ( .B1(n260), .B2(n297), .C1(n298), .C2(n265), .A(n299), .ZN(
        n296) );
  INV_X1 U464 ( .A(n305), .ZN(n297) );
  NAND2_X1 U465 ( .A1(n452), .A2(n453), .ZN(OUTSHFT[21]) );
  AOI221_X1 U466 ( .B1(n627), .B2(n206), .C1(n243), .C2(n211), .A(n461), .ZN(
        n452) );
  AOI221_X1 U467 ( .B1(n258), .B2(n210), .C1(n205), .C2(n265), .A(n454), .ZN(
        n453) );
  OAI22_X1 U468 ( .A1(n202), .A2(n462), .B1(n463), .B2(n329), .ZN(n461) );
  INV_X1 U469 ( .A(n465), .ZN(n202) );
  OAI221_X1 U470 ( .B1(n363), .B2(n290), .C1(n356), .C2(n124), .A(n466), .ZN(
        n465) );
  AOI22_X1 U471 ( .A1(n134), .A2(n366), .B1(n597), .B2(n467), .ZN(n466) );
  OR3_X1 U472 ( .A1(n175), .A2(n737), .A3(n319), .ZN(n654) );
  INV_X1 U473 ( .A(n232), .ZN(n231) );
  AOI22_X1 U474 ( .A1(n233), .A2(n234), .B1(n235), .B2(n236), .ZN(n232) );
  INV_X1 U475 ( .A(n491), .ZN(n490) );
  AOI22_X1 U476 ( .A1(n492), .A2(n229), .B1(n493), .B2(n227), .ZN(n491) );
  INV_X1 U477 ( .A(n275), .ZN(n274) );
  AOI22_X1 U478 ( .A1(n276), .A2(n229), .B1(n277), .B2(n227), .ZN(n275) );
  BUF_X1 U479 ( .A(n342), .Z(n587) );
  BUF_X1 U480 ( .A(n342), .Z(n557) );
  BUF_X1 U481 ( .A(n342), .Z(n585) );
  INV_X1 U482 ( .A(n590), .ZN(n109) );
  OAI22_X1 U483 ( .A1(n600), .A2(n112), .B1(n601), .B2(n106), .ZN(n599) );
  OAI22_X1 U484 ( .A1(n595), .A2(n584), .B1(n621), .B2(n117), .ZN(n695) );
  OAI22_X1 U485 ( .A1(n619), .A2(n113), .B1(n664), .B2(n105), .ZN(n663) );
  OAI22_X1 U486 ( .A1(n97), .A2(n112), .B1(n96), .B2(n105), .ZN(n615) );
  OAI22_X1 U487 ( .A1(n89), .A2(n114), .B1(n669), .B2(n106), .ZN(n705) );
  OAI22_X1 U488 ( .A1(n621), .A2(n113), .B1(n107), .B2(n673), .ZN(n718) );
  OAI22_X1 U489 ( .A1(n623), .A2(n112), .B1(n592), .B2(n107), .ZN(n726) );
  NAND2_X1 U490 ( .A1(n301), .A2(n329), .ZN(n162) );
  OAI221_X1 U491 ( .B1(n119), .B2(n719), .C1(n117), .C2(n101), .A(n682), .ZN(
        n235) );
  OAI221_X1 U492 ( .B1(n120), .B2(n100), .C1(n117), .C2(n99), .A(n632), .ZN(
        n366) );
  AOI221_X1 U493 ( .B1(n121), .B2(DATA1[29]), .C1(DATA1[28]), .C2(n118), .A(
        n701), .ZN(n574) );
  OAI22_X1 U494 ( .A1(n664), .A2(n114), .B1(n619), .B2(n107), .ZN(n701) );
  OAI221_X1 U495 ( .B1(n584), .B2(n592), .C1(n586), .C2(n591), .A(n716), .ZN(
        n382) );
  AOI22_X1 U496 ( .A1(DATA1[16]), .A2(n110), .B1(DATA1[17]), .B2(n104), .ZN(
        n716) );
  OAI221_X1 U497 ( .B1(n584), .B2(n89), .C1(n586), .C2(n90), .A(n677), .ZN(
        n421) );
  AOI22_X1 U498 ( .A1(DATA1[11]), .A2(n111), .B1(DATA1[12]), .B2(n103), .ZN(
        n677) );
  OAI221_X1 U499 ( .B1(n119), .B2(n90), .C1(n586), .C2(n89), .A(n734), .ZN(
        n387) );
  AOI22_X1 U500 ( .A1(DATA1[16]), .A2(n110), .B1(DATA1[15]), .B2(n103), .ZN(
        n734) );
  OAI221_X1 U501 ( .B1(n120), .B2(n595), .C1(n586), .C2(n594), .A(n715), .ZN(
        n383) );
  AOI22_X1 U502 ( .A1(DATA1[20]), .A2(n111), .B1(DATA1[21]), .B2(n104), .ZN(
        n715) );
  OAI221_X1 U503 ( .B1(n584), .B2(n98), .C1(n586), .C2(n99), .A(n608), .ZN(
        n370) );
  OAI221_X1 U504 ( .B1(n120), .B2(n97), .C1(n117), .C2(n98), .A(n697), .ZN(
        n439) );
  AOI21_X1 U505 ( .B1(DATA1[3]), .B2(n104), .A(n698), .ZN(n697) );
  OAI221_X1 U506 ( .B1(n119), .B2(n661), .C1(n117), .C2(n623), .A(n704), .ZN(
        n443) );
  AOI22_X1 U507 ( .A1(DATA1[18]), .A2(n110), .B1(DATA1[19]), .B2(n103), .ZN(
        n704) );
  OAI221_X1 U508 ( .B1(n119), .B2(n619), .C1(n601), .C2(n117), .A(n710), .ZN(
        n448) );
  AOI21_X1 U509 ( .B1(DATA1[29]), .B2(n104), .A(n689), .ZN(n710) );
  OAI221_X1 U510 ( .B1(n584), .B2(n594), .C1(n586), .C2(n661), .A(n675), .ZN(
        n420) );
  AOI22_X1 U511 ( .A1(DATA1[19]), .A2(n111), .B1(DATA1[20]), .B2(n103), .ZN(
        n675) );
  AOI211_X1 U512 ( .C1(n121), .C2(DATA1[1]), .A(n699), .B(n688), .ZN(n436) );
  OAI221_X1 U513 ( .B1(n120), .B2(n611), .C1(n117), .C2(n600), .A(n667), .ZN(
        n415) );
  AOI22_X1 U514 ( .A1(DATA1[27]), .A2(n111), .B1(DATA1[28]), .B2(n590), .ZN(
        n667) );
  OAI221_X1 U515 ( .B1(n584), .B2(n92), .C1(n117), .C2(n91), .A(n692), .ZN(
        n433) );
  OAI221_X1 U516 ( .B1(n120), .B2(n601), .C1(n117), .C2(n600), .A(n683), .ZN(
        n403) );
  AOI21_X1 U517 ( .B1(DATA1[30]), .B2(n103), .A(n655), .ZN(n683) );
  OAI221_X1 U518 ( .B1(n673), .B2(n584), .C1(n117), .C2(n621), .A(n703), .ZN(
        n451) );
  AOI22_X1 U519 ( .A1(DATA1[22]), .A2(n111), .B1(DATA1[23]), .B2(n103), .ZN(
        n703) );
  OAI221_X1 U520 ( .B1(n664), .B2(n119), .C1(n673), .C2(n586), .A(n674), .ZN(
        n416) );
  AOI22_X1 U521 ( .A1(DATA1[23]), .A2(n111), .B1(DATA1[24]), .B2(n590), .ZN(
        n674) );
  OAI221_X1 U522 ( .B1(n120), .B2(n601), .C1(n586), .C2(n619), .A(n620), .ZN(
        n371) );
  AOI22_X1 U523 ( .A1(DATA1[25]), .A2(n110), .B1(DATA1[26]), .B2(n590), .ZN(
        n620) );
  OAI221_X1 U524 ( .B1(n119), .B2(n96), .C1(n117), .C2(n95), .A(n628), .ZN(
        n365) );
  AOI22_X1 U525 ( .A1(DATA1[9]), .A2(n110), .B1(DATA1[8]), .B2(n590), .ZN(n628) );
  OAI221_X1 U526 ( .B1(n584), .B2(n621), .C1(n117), .C2(n595), .A(n622), .ZN(
        n353) );
  AOI22_X1 U527 ( .A1(DATA1[21]), .A2(n110), .B1(DATA1[22]), .B2(n104), .ZN(
        n622) );
  OAI221_X1 U528 ( .B1(n119), .B2(n99), .C1(n586), .C2(n98), .A(n708), .ZN(
        n449) );
  OAI221_X1 U529 ( .B1(n584), .B2(n101), .C1(n586), .C2(n100), .A(n731), .ZN(
        n392) );
  AOI22_X1 U530 ( .A1(DATA1[4]), .A2(n111), .B1(DATA1[3]), .B2(n104), .ZN(n731) );
  INV_X1 U531 ( .A(n339), .ZN(n173) );
  INV_X1 U532 ( .A(n301), .ZN(n243) );
  OAI221_X1 U533 ( .B1(n119), .B2(n625), .C1(n586), .C2(n659), .A(n660), .ZN(
        n410) );
  AOI22_X1 U534 ( .A1(DATA1[19]), .A2(n111), .B1(DATA1[18]), .B2(n590), .ZN(
        n660) );
  OAI221_X1 U535 ( .B1(n120), .B2(n591), .C1(n586), .C2(n592), .A(n593), .ZN(
        n360) );
  AOI22_X1 U536 ( .A1(DATA1[21]), .A2(n110), .B1(DATA1[20]), .B2(n104), .ZN(
        n593) );
  OAI221_X1 U537 ( .B1(n584), .B2(n669), .C1(n117), .C2(n625), .A(n693), .ZN(
        n432) );
  AOI22_X1 U538 ( .A1(DATA1[18]), .A2(n110), .B1(DATA1[17]), .B2(n103), .ZN(
        n693) );
  OAI221_X1 U539 ( .B1(n119), .B2(n669), .C1(n586), .C2(n89), .A(n721), .ZN(
        n482) );
  OAI221_X1 U540 ( .B1(n119), .B2(n625), .C1(n117), .C2(n669), .A(n626), .ZN(
        n355) );
  OAI221_X1 U541 ( .B1(n584), .B2(n91), .C1(n117), .C2(n90), .A(n658), .ZN(
        n411) );
  AOI22_X1 U542 ( .A1(DATA1[15]), .A2(n110), .B1(DATA1[14]), .B2(n590), .ZN(
        n658) );
  OAI221_X1 U543 ( .B1(n120), .B2(n89), .C1(n117), .C2(n669), .A(n588), .ZN(
        n362) );
  AOI22_X1 U544 ( .A1(DATA1[17]), .A2(n111), .B1(DATA1[16]), .B2(n103), .ZN(
        n588) );
  OAI221_X1 U545 ( .B1(n120), .B2(n94), .C1(n586), .C2(n93), .A(n733), .ZN(
        n388) );
  AOI22_X1 U546 ( .A1(DATA1[12]), .A2(n111), .B1(DATA1[11]), .B2(n104), .ZN(
        n733) );
  OAI221_X1 U547 ( .B1(n120), .B2(n661), .C1(n586), .C2(n594), .A(n727), .ZN(
        n478) );
  AOI22_X1 U548 ( .A1(DATA1[24]), .A2(n110), .B1(DATA1[23]), .B2(n104), .ZN(
        n727) );
  OAI221_X1 U549 ( .B1(n584), .B2(n93), .C1(n117), .C2(n92), .A(n630), .ZN(
        n460) );
  OAI221_X1 U550 ( .B1(n119), .B2(n97), .C1(n586), .C2(n96), .A(n732), .ZN(
        n393) );
  AOI22_X1 U551 ( .A1(DATA1[8]), .A2(n110), .B1(DATA1[7]), .B2(n104), .ZN(n732) );
  OAI221_X1 U552 ( .B1(n120), .B2(n623), .C1(n586), .C2(n592), .A(n624), .ZN(
        n471) );
  AOI22_X1 U553 ( .A1(DATA1[17]), .A2(n110), .B1(DATA1[18]), .B2(n590), .ZN(
        n624) );
  OAI22_X1 U554 ( .A1(n655), .A2(n641), .B1(DATA2[2]), .B2(n415), .ZN(n319) );
  OAI221_X1 U555 ( .B1(n584), .B2(n246), .C1(n586), .C2(n611), .A(n717), .ZN(
        n303) );
  AOI22_X1 U556 ( .A1(DATA1[28]), .A2(n111), .B1(DATA1[29]), .B2(n104), .ZN(
        n717) );
  AOI21_X1 U557 ( .B1(DATA2[1]), .B2(n102), .A(n604), .ZN(n341) );
  OAI221_X1 U558 ( .B1(n584), .B2(n594), .C1(n586), .C2(n595), .A(n596), .ZN(
        n542) );
  AOI22_X1 U559 ( .A1(DATA1[25]), .A2(n110), .B1(DATA1[24]), .B2(n104), .ZN(
        n596) );
  OAI221_X1 U560 ( .B1(n120), .B2(n623), .C1(n586), .C2(n661), .A(n662), .ZN(
        n559) );
  AOI22_X1 U561 ( .A1(DATA1[23]), .A2(n111), .B1(DATA1[22]), .B2(n590), .ZN(
        n662) );
  OAI221_X1 U562 ( .B1(n119), .B2(n680), .C1(n117), .C2(n94), .A(n681), .ZN(
        n511) );
  AOI22_X1 U563 ( .A1(DATA1[11]), .A2(n111), .B1(DATA1[10]), .B2(n103), .ZN(
        n681) );
  OAI221_X1 U564 ( .B1(n119), .B2(n592), .C1(n117), .C2(n623), .A(n694), .ZN(
        n570) );
  AOI22_X1 U565 ( .A1(DATA1[22]), .A2(n110), .B1(DATA1[21]), .B2(n103), .ZN(
        n694) );
  OAI221_X1 U566 ( .B1(n120), .B2(n92), .C1(n117), .C2(n93), .A(n722), .ZN(
        n643) );
  AOI22_X1 U567 ( .A1(DATA1[8]), .A2(n110), .B1(DATA1[9]), .B2(n104), .ZN(n722) );
  OAI221_X1 U568 ( .B1(n119), .B2(n90), .C1(n117), .C2(n91), .A(n706), .ZN(
        n444) );
  AOI22_X1 U569 ( .A1(DATA1[10]), .A2(n111), .B1(DATA1[11]), .B2(n103), .ZN(
        n706) );
  OAI221_X1 U570 ( .B1(n120), .B2(n591), .C1(n117), .C2(n659), .A(n676), .ZN(
        n518) );
  AOI22_X1 U571 ( .A1(DATA1[15]), .A2(n111), .B1(DATA1[16]), .B2(n590), .ZN(
        n676) );
  OAI221_X1 U572 ( .B1(n673), .B2(n120), .C1(n664), .C2(n586), .A(n728), .ZN(
        n650) );
  AOI22_X1 U573 ( .A1(DATA1[28]), .A2(n111), .B1(DATA1[27]), .B2(n104), .ZN(
        n728) );
  OAI22_X1 U574 ( .A1(n641), .A2(n377), .B1(DATA2[2]), .B2(n642), .ZN(n221) );
  NAND2_X1 U575 ( .A1(n250), .A2(n254), .ZN(n186) );
  NAND2_X1 U576 ( .A1(DATA2[4]), .A2(n497), .ZN(n175) );
  NAND2_X1 U577 ( .A1(n160), .A2(n498), .ZN(n197) );
  OAI22_X1 U578 ( .A1(n213), .A2(n462), .B1(n476), .B2(n301), .ZN(n475) );
  INV_X1 U579 ( .A(n223), .ZN(n476) );
  INV_X1 U580 ( .A(DATA2[4]), .ZN(n254) );
  NAND2_X1 U581 ( .A1(n251), .A2(DATA2[4]), .ZN(n462) );
  INV_X1 U582 ( .A(DATA1[30]), .ZN(n611) );
  NAND2_X1 U583 ( .A1(DATA2[1]), .A2(n736), .ZN(n586) );
  NAND2_X1 U584 ( .A1(n301), .A2(n495), .ZN(n234) );
  OAI21_X1 U585 ( .B1(n496), .B2(n494), .A(n254), .ZN(n495) );
  INV_X1 U586 ( .A(n245), .ZN(n496) );
  NOR2_X1 U587 ( .A1(n736), .A2(DATA2[1]), .ZN(n590) );
  INV_X1 U588 ( .A(DATA1[29]), .ZN(n600) );
  INV_X1 U589 ( .A(DATA1[19]), .ZN(n592) );
  INV_X1 U590 ( .A(DATA1[20]), .ZN(n623) );
  OAI21_X1 U591 ( .B1(n300), .B2(n301), .A(n302), .ZN(n299) );
  INV_X1 U592 ( .A(n304), .ZN(n300) );
  NAND2_X1 U593 ( .A1(n497), .A2(n254), .ZN(n329) );
  OAI211_X1 U594 ( .C1(n551), .C2(n552), .A(n553), .B(n554), .ZN(OUTSHFT[15])
         );
  INV_X1 U595 ( .A(n242), .ZN(n551) );
  AOI22_X1 U596 ( .A1(n253), .A2(n265), .B1(n241), .B2(n162), .ZN(n553) );
  AOI211_X1 U597 ( .C1(n634), .C2(n252), .A(n339), .B(n555), .ZN(n554) );
  NAND2_X1 U598 ( .A1(n289), .A2(n498), .ZN(n314) );
  INV_X1 U599 ( .A(DATA2[2]), .ZN(n641) );
  INV_X1 U600 ( .A(DATA1[26]), .ZN(n664) );
  INV_X1 U601 ( .A(DATA1[22]), .ZN(n594) );
  INV_X1 U602 ( .A(DATA1[25]), .ZN(n673) );
  INV_X1 U603 ( .A(DATA1[23]), .ZN(n595) );
  INV_X1 U604 ( .A(DATA1[27]), .ZN(n619) );
  INV_X1 U605 ( .A(DATA1[21]), .ZN(n661) );
  INV_X1 U606 ( .A(DATA1[24]), .ZN(n621) );
  INV_X1 U607 ( .A(DATA1[28]), .ZN(n601) );
  INV_X1 U623 ( .A(DATA1[18]), .ZN(n591) );
  INV_X1 U624 ( .A(n552), .ZN(n163) );
  INV_X1 U625 ( .A(DATA1[16]), .ZN(n625) );
  NAND2_X1 U626 ( .A1(n497), .A2(n498), .ZN(n245) );
  NAND2_X1 U627 ( .A1(n250), .A2(DATA2[4]), .ZN(n455) );
  AND2_X1 U628 ( .A1(n494), .A2(DATA2[4]), .ZN(n229) );
  NAND2_X1 U629 ( .A1(n737), .A2(DATA2[2]), .ZN(n358) );
  NAND2_X1 U630 ( .A1(DATA2[2]), .A2(n738), .ZN(n342) );
  NAND2_X1 U631 ( .A1(n552), .A2(n175), .ZN(n644) );
  AOI22_X1 U632 ( .A1(n243), .A2(n164), .B1(n657), .B2(n165), .ZN(n335) );
  AOI22_X1 U633 ( .A1(n154), .A2(n265), .B1(n629), .B2(n161), .ZN(n336) );
  AOI211_X1 U634 ( .C1(n289), .C2(n159), .A(n338), .B(n339), .ZN(n337) );
  INV_X1 U635 ( .A(DATA1[17]), .ZN(n659) );
  NAND2_X1 U636 ( .A1(DATA2[1]), .A2(n735), .ZN(n584) );
  INV_X1 U637 ( .A(DATA2[3]), .ZN(n738) );
  OAI22_X1 U638 ( .A1(n99), .A2(n114), .B1(n98), .B2(n106), .ZN(n670) );
  OR2_X1 U639 ( .A1(n713), .A2(n711), .ZN(n724) );
  INV_X1 U640 ( .A(n240), .ZN(OUTSHFT[31]) );
  AOI221_X1 U641 ( .B1(n241), .B2(n629), .C1(n242), .C2(n243), .A(n244), .ZN(
        n240) );
  OAI221_X1 U642 ( .B1(n245), .B2(n246), .C1(n247), .C2(n248), .A(n249), .ZN(
        n244) );
  OAI222_X1 U643 ( .A1(n250), .A2(n251), .B1(n252), .B2(DATA2[4]), .C1(n253), 
        .C2(n254), .ZN(n249) );
  OR2_X1 U644 ( .A1(DATA2[1]), .A2(n735), .ZN(n88) );
  BUF_X1 U645 ( .A(DATA1[31]), .Z(n102) );
  NOR2_X1 U646 ( .A1(n739), .A2(FUNC[1]), .ZN(n497) );
  NOR2_X1 U647 ( .A1(n556), .A2(US), .ZN(n339) );
  NOR2_X1 U648 ( .A1(FUNC[0]), .A2(FUNC[1]), .ZN(n250) );
  AND2_X1 U649 ( .A1(FUNC[1]), .A2(n739), .ZN(n251) );
  INV_X1 U650 ( .A(US), .ZN(n498) );
  OAI211_X1 U651 ( .C1(n635), .C2(n462), .A(n636), .B(n637), .ZN(OUTSHFT[12])
         );
  AND2_X1 U652 ( .A1(US), .A2(n497), .ZN(n494) );
  INV_X1 U653 ( .A(DATA1[14]), .ZN(n89) );
  INV_X1 U654 ( .A(DATA1[13]), .ZN(n90) );
  INV_X1 U655 ( .A(DATA1[12]), .ZN(n91) );
  INV_X1 U656 ( .A(DATA1[11]), .ZN(n92) );
  INV_X1 U657 ( .A(DATA1[10]), .ZN(n93) );
  INV_X1 U658 ( .A(DATA1[9]), .ZN(n94) );
  INV_X1 U659 ( .A(DATA1[7]), .ZN(n95) );
  INV_X1 U660 ( .A(DATA1[6]), .ZN(n96) );
  INV_X1 U661 ( .A(DATA1[5]), .ZN(n97) );
  INV_X1 U662 ( .A(DATA1[4]), .ZN(n98) );
  INV_X1 U663 ( .A(DATA1[3]), .ZN(n99) );
  INV_X1 U664 ( .A(DATA1[2]), .ZN(n100) );
  INV_X1 U665 ( .A(DATA1[1]), .ZN(n101) );
  INV_X1 U666 ( .A(DATA2[0]), .ZN(n736) );
  AOI22_X1 U667 ( .A1(DATA1[12]), .A2(n110), .B1(DATA1[13]), .B2(n104), .ZN(
        n721) );
  AOI22_X1 U668 ( .A1(DATA1[14]), .A2(n111), .B1(DATA1[13]), .B2(n103), .ZN(
        n692) );
  AOI22_X1 U669 ( .A1(DATA1[13]), .A2(n110), .B1(DATA1[14]), .B2(n103), .ZN(
        n626) );
  AOI22_X1 U670 ( .A1(DATA1[13]), .A2(n110), .B1(DATA1[12]), .B2(n590), .ZN(
        n630) );
  AOI22_X1 U671 ( .A1(DATA1[3]), .A2(n111), .B1(DATA1[2]), .B2(n103), .ZN(n682) );
  AOI21_X1 U672 ( .B1(DATA1[2]), .B2(n104), .A(n609), .ZN(n608) );
  AOI22_X1 U673 ( .A1(DATA1[6]), .A2(n110), .B1(DATA1[5]), .B2(n104), .ZN(n708) );
  AOI22_X1 U674 ( .A1(DATA1[5]), .A2(n110), .B1(DATA1[4]), .B2(n104), .ZN(n632) );
  NAND2_X1 U675 ( .A1(DATA1[0]), .A2(n111), .ZN(n377) );
  CLKBUF_X1 U676 ( .A(n584), .Z(n119) );
  CLKBUF_X1 U677 ( .A(n584), .Z(n120) );
  INV_X1 U678 ( .A(n120), .ZN(n121) );
  INV_X1 U679 ( .A(n122), .ZN(n126) );
  INV_X1 U680 ( .A(n123), .ZN(n127) );
  INV_X1 U681 ( .A(DATA1[15]), .ZN(n669) );
  INV_X1 U682 ( .A(DATA1[8]), .ZN(n680) );
  INV_X1 U683 ( .A(DATA1[0]), .ZN(n719) );
  INV_X1 U684 ( .A(n736), .ZN(n735) );
  INV_X1 U685 ( .A(n738), .ZN(n737) );
  INV_X1 U686 ( .A(FUNC[0]), .ZN(n739) );
endmodule


module BOOTHMUL_NB32 ( A, B, C );
  input [15:0] A;
  input [15:0] B;
  output [31:0] C;
  wire   \Term[7][31] , \Term[7][30] , \Term[7][29] , \Term[7][28] ,
         \Term[7][27] , \Term[7][26] , \Term[7][25] , \Term[7][24] ,
         \Term[7][23] , \Term[7][22] , \Term[7][21] , \Term[7][20] ,
         \Term[7][19] , \Term[7][18] , \Term[7][17] , \Term[7][16] ,
         \Term[7][15] , \Term[7][14] , \Term[7][13] , \Term[7][12] ,
         \Term[7][11] , \Term[7][10] , \Term[7][9] , \Term[7][8] ,
         \Term[7][7] , \Term[7][6] , \Term[7][5] , \Term[7][4] , \Term[7][3] ,
         \Term[7][2] , \Term[7][1] , \Term[7][0] , \Term[6][31] ,
         \Term[6][30] , \Term[6][29] , \Term[6][28] , \Term[6][27] ,
         \Term[6][26] , \Term[6][25] , \Term[6][24] , \Term[6][23] ,
         \Term[6][22] , \Term[6][21] , \Term[6][20] , \Term[6][19] ,
         \Term[6][18] , \Term[6][17] , \Term[6][16] , \Term[6][15] ,
         \Term[6][14] , \Term[6][13] , \Term[6][12] , \Term[6][11] ,
         \Term[6][10] , \Term[6][9] , \Term[6][8] , \Term[6][7] , \Term[6][6] ,
         \Term[6][5] , \Term[6][4] , \Term[6][3] , \Term[6][2] , \Term[6][1] ,
         \Term[6][0] , \Term[5][31] , \Term[5][30] , \Term[5][29] ,
         \Term[5][28] , \Term[5][27] , \Term[5][26] , \Term[5][25] ,
         \Term[5][24] , \Term[5][23] , \Term[5][22] , \Term[5][21] ,
         \Term[5][20] , \Term[5][19] , \Term[5][18] , \Term[5][17] ,
         \Term[5][16] , \Term[5][15] , \Term[5][14] , \Term[5][13] ,
         \Term[5][12] , \Term[5][11] , \Term[5][10] , \Term[5][9] ,
         \Term[5][8] , \Term[5][7] , \Term[5][6] , \Term[5][5] , \Term[5][4] ,
         \Term[5][3] , \Term[5][2] , \Term[5][1] , \Term[5][0] , \Term[4][31] ,
         \Term[4][30] , \Term[4][29] , \Term[4][28] , \Term[4][27] ,
         \Term[4][26] , \Term[4][25] , \Term[4][24] , \Term[4][23] ,
         \Term[4][22] , \Term[4][21] , \Term[4][20] , \Term[4][19] ,
         \Term[4][18] , \Term[4][17] , \Term[4][16] , \Term[4][15] ,
         \Term[4][14] , \Term[4][13] , \Term[4][12] , \Term[4][11] ,
         \Term[4][10] , \Term[4][9] , \Term[4][8] , \Term[4][7] , \Term[4][6] ,
         \Term[4][5] , \Term[4][4] , \Term[4][3] , \Term[4][2] , \Term[4][1] ,
         \Term[4][0] , \Term[3][31] , \Term[3][30] , \Term[3][29] ,
         \Term[3][28] , \Term[3][27] , \Term[3][26] , \Term[3][25] ,
         \Term[3][24] , \Term[3][23] , \Term[3][22] , \Term[3][21] ,
         \Term[3][20] , \Term[3][19] , \Term[3][18] , \Term[3][17] ,
         \Term[3][16] , \Term[3][15] , \Term[3][14] , \Term[3][13] ,
         \Term[3][12] , \Term[3][11] , \Term[3][10] , \Term[3][9] ,
         \Term[3][8] , \Term[3][7] , \Term[3][6] , \Term[3][5] , \Term[3][4] ,
         \Term[3][3] , \Term[3][2] , \Term[3][1] , \Term[3][0] , \Term[2][31] ,
         \Term[2][30] , \Term[2][29] , \Term[2][28] , \Term[2][27] ,
         \Term[2][26] , \Term[2][25] , \Term[2][24] , \Term[2][23] ,
         \Term[2][22] , \Term[2][21] , \Term[2][20] , \Term[2][19] ,
         \Term[2][18] , \Term[2][17] , \Term[2][16] , \Term[2][15] ,
         \Term[2][14] , \Term[2][13] , \Term[2][12] , \Term[2][11] ,
         \Term[2][10] , \Term[2][9] , \Term[2][8] , \Term[2][7] , \Term[2][6] ,
         \Term[2][5] , \Term[2][4] , \Term[2][3] , \Term[2][2] , \Term[2][1] ,
         \Term[2][0] , \Term[1][31] , \Term[1][30] , \Term[1][29] ,
         \Term[1][28] , \Term[1][27] , \Term[1][26] , \Term[1][25] ,
         \Term[1][24] , \Term[1][23] , \Term[1][22] , \Term[1][21] ,
         \Term[1][20] , \Term[1][19] , \Term[1][18] , \Term[1][17] ,
         \Term[1][16] , \Term[1][15] , \Term[1][14] , \Term[1][13] ,
         \Term[1][12] , \Term[1][11] , \Term[1][10] , \Term[1][9] ,
         \Term[1][8] , \Term[1][7] , \Term[1][6] , \Term[1][5] , \Term[1][4] ,
         \Term[1][3] , \Term[1][2] , \Term[1][1] , \Term[1][0] , \Term[0][31] ,
         \Term[0][30] , \Term[0][29] , \Term[0][28] , \Term[0][27] ,
         \Term[0][26] , \Term[0][25] , \Term[0][24] , \Term[0][23] ,
         \Term[0][22] , \Term[0][21] , \Term[0][20] , \Term[0][19] ,
         \Term[0][18] , \Term[0][17] , \Term[0][16] , \Term[0][15] ,
         \Term[0][14] , \Term[0][13] , \Term[0][12] , \Term[0][11] ,
         \Term[0][10] , \Term[0][9] , \Term[0][8] , \Term[0][7] , \Term[0][6] ,
         \Term[0][5] , \Term[0][4] , \Term[0][3] , \Term[0][2] , \Term[0][1] ,
         \Term[0][0] , \Res[6][31] , \Res[6][30] , \Res[6][29] , \Res[6][28] ,
         \Res[6][27] , \Res[6][26] , \Res[6][25] , \Res[6][24] , \Res[6][23] ,
         \Res[6][22] , \Res[6][21] , \Res[6][20] , \Res[6][19] , \Res[6][18] ,
         \Res[6][17] , \Res[6][16] , \Res[6][15] , \Res[6][14] , \Res[6][13] ,
         \Res[6][12] , \Res[6][11] , \Res[6][10] , \Res[6][9] , \Res[6][8] ,
         \Res[6][7] , \Res[6][6] , \Res[6][5] , \Res[6][4] , \Res[6][3] ,
         \Res[6][2] , \Res[6][1] , \Res[6][0] , \Res[5][31] , \Res[5][30] ,
         \Res[5][29] , \Res[5][28] , \Res[5][27] , \Res[5][26] , \Res[5][25] ,
         \Res[5][24] , \Res[5][23] , \Res[5][22] , \Res[5][21] , \Res[5][20] ,
         \Res[5][19] , \Res[5][18] , \Res[5][17] , \Res[5][16] , \Res[5][15] ,
         \Res[5][14] , \Res[5][13] , \Res[5][12] , \Res[5][11] , \Res[5][10] ,
         \Res[5][9] , \Res[5][8] , \Res[5][7] , \Res[5][6] , \Res[5][5] ,
         \Res[5][4] , \Res[5][3] , \Res[5][2] , \Res[5][1] , \Res[5][0] ,
         \Res[4][31] , \Res[4][30] , \Res[4][29] , \Res[4][28] , \Res[4][27] ,
         \Res[4][26] , \Res[4][25] , \Res[4][24] , \Res[4][23] , \Res[4][22] ,
         \Res[4][21] , \Res[4][20] , \Res[4][19] , \Res[4][18] , \Res[4][17] ,
         \Res[4][16] , \Res[4][15] , \Res[4][14] , \Res[4][13] , \Res[4][12] ,
         \Res[4][11] , \Res[4][10] , \Res[4][9] , \Res[4][8] , \Res[4][7] ,
         \Res[4][6] , \Res[4][5] , \Res[4][4] , \Res[4][3] , \Res[4][2] ,
         \Res[4][1] , \Res[4][0] , \Res[3][31] , \Res[3][30] , \Res[3][29] ,
         \Res[3][28] , \Res[3][27] , \Res[3][26] , \Res[3][25] , \Res[3][24] ,
         \Res[3][23] , \Res[3][22] , \Res[3][21] , \Res[3][20] , \Res[3][19] ,
         \Res[3][18] , \Res[3][17] , \Res[3][16] , \Res[3][15] , \Res[3][14] ,
         \Res[3][13] , \Res[3][12] , \Res[3][11] , \Res[3][10] , \Res[3][9] ,
         \Res[3][8] , \Res[3][7] , \Res[3][6] , \Res[3][5] , \Res[3][4] ,
         \Res[3][3] , \Res[3][2] , \Res[3][1] , \Res[3][0] , \Res[2][31] ,
         \Res[2][30] , \Res[2][29] , \Res[2][28] , \Res[2][27] , \Res[2][26] ,
         \Res[2][25] , \Res[2][24] , \Res[2][23] , \Res[2][22] , \Res[2][21] ,
         \Res[2][20] , \Res[2][19] , \Res[2][18] , \Res[2][17] , \Res[2][16] ,
         \Res[2][15] , \Res[2][14] , \Res[2][13] , \Res[2][12] , \Res[2][11] ,
         \Res[2][10] , \Res[2][9] , \Res[2][8] , \Res[2][7] , \Res[2][6] ,
         \Res[2][5] , \Res[2][4] , \Res[2][3] , \Res[2][2] , \Res[2][1] ,
         \Res[2][0] , \Res[1][31] , \Res[1][30] , \Res[1][29] , \Res[1][28] ,
         \Res[1][27] , \Res[1][26] , \Res[1][25] , \Res[1][24] , \Res[1][23] ,
         \Res[1][22] , \Res[1][21] , \Res[1][20] , \Res[1][19] , \Res[1][18] ,
         \Res[1][17] , \Res[1][16] , \Res[1][15] , \Res[1][14] , \Res[1][13] ,
         \Res[1][12] , \Res[1][11] , \Res[1][10] , \Res[1][9] , \Res[1][8] ,
         \Res[1][7] , \Res[1][6] , \Res[1][5] , \Res[1][4] , \Res[1][3] ,
         \Res[1][2] , \Res[1][1] , \Res[1][0] , \Res[0][31] , \Res[0][30] ,
         \Res[0][29] , \Res[0][28] , \Res[0][27] , \Res[0][26] , \Res[0][25] ,
         \Res[0][24] , \Res[0][23] , \Res[0][22] , \Res[0][21] , \Res[0][20] ,
         \Res[0][19] , \Res[0][18] , \Res[0][17] , \Res[0][16] , \Res[0][15] ,
         \Res[0][14] , \Res[0][13] , \Res[0][12] , \Res[0][11] , \Res[0][10] ,
         \Res[0][9] , \Res[0][8] , \Res[0][7] , \Res[0][6] , \Res[0][5] ,
         \Res[0][4] , \Res[0][3] , \Res[0][2] , \Res[0][1] , \Res[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] OP;
  assign n1 = A[0];
  assign n2 = A[1];
  assign n3 = A[2];
  assign n4 = A[3];
  assign n5 = A[4];
  assign n6 = A[5];
  assign n7 = A[6];
  assign n8 = A[7];
  assign n9 = A[8];
  assign n10 = A[9];
  assign n11 = A[10];
  assign n12 = A[11];
  assign n13 = A[12];
  assign n14 = A[13];
  assign n15 = A[14];

  MUX_SHIFT_NB16_N_sh0 mux_map_0 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel({B[1:0], 1'b0}), .AS(OP[0]), 
        .B({\Term[0][31] , \Term[0][30] , \Term[0][29] , \Term[0][28] , 
        \Term[0][27] , \Term[0][26] , \Term[0][25] , \Term[0][24] , 
        \Term[0][23] , \Term[0][22] , \Term[0][21] , \Term[0][20] , 
        \Term[0][19] , \Term[0][18] , \Term[0][17] , \Term[0][16] , 
        \Term[0][15] , \Term[0][14] , \Term[0][13] , \Term[0][12] , 
        \Term[0][11] , \Term[0][10] , \Term[0][9] , \Term[0][8] , \Term[0][7] , 
        \Term[0][6] , \Term[0][5] , \Term[0][4] , \Term[0][3] , \Term[0][2] , 
        \Term[0][1] , \Term[0][0] }) );
  MUX_SHIFT_NB16_N_sh2 mux_map_1 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel(B[3:1]), .AS(OP[1]), .B({
        \Term[1][31] , \Term[1][30] , \Term[1][29] , \Term[1][28] , 
        \Term[1][27] , \Term[1][26] , \Term[1][25] , \Term[1][24] , 
        \Term[1][23] , \Term[1][22] , \Term[1][21] , \Term[1][20] , 
        \Term[1][19] , \Term[1][18] , \Term[1][17] , \Term[1][16] , 
        \Term[1][15] , \Term[1][14] , \Term[1][13] , \Term[1][12] , 
        \Term[1][11] , \Term[1][10] , \Term[1][9] , \Term[1][8] , \Term[1][7] , 
        \Term[1][6] , \Term[1][5] , \Term[1][4] , \Term[1][3] , \Term[1][2] , 
        \Term[1][1] , \Term[1][0] }) );
  MUX_SHIFT_NB16_N_sh4 mux_map_2 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel(B[5:3]), .AS(OP[2]), .B({
        \Term[2][31] , \Term[2][30] , \Term[2][29] , \Term[2][28] , 
        \Term[2][27] , \Term[2][26] , \Term[2][25] , \Term[2][24] , 
        \Term[2][23] , \Term[2][22] , \Term[2][21] , \Term[2][20] , 
        \Term[2][19] , \Term[2][18] , \Term[2][17] , \Term[2][16] , 
        \Term[2][15] , \Term[2][14] , \Term[2][13] , \Term[2][12] , 
        \Term[2][11] , \Term[2][10] , \Term[2][9] , \Term[2][8] , \Term[2][7] , 
        \Term[2][6] , \Term[2][5] , \Term[2][4] , \Term[2][3] , \Term[2][2] , 
        \Term[2][1] , \Term[2][0] }) );
  MUX_SHIFT_NB16_N_sh6 mux_map_3 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel(B[7:5]), .AS(OP[3]), .B({
        \Term[3][31] , \Term[3][30] , \Term[3][29] , \Term[3][28] , 
        \Term[3][27] , \Term[3][26] , \Term[3][25] , \Term[3][24] , 
        \Term[3][23] , \Term[3][22] , \Term[3][21] , \Term[3][20] , 
        \Term[3][19] , \Term[3][18] , \Term[3][17] , \Term[3][16] , 
        \Term[3][15] , \Term[3][14] , \Term[3][13] , \Term[3][12] , 
        \Term[3][11] , \Term[3][10] , \Term[3][9] , \Term[3][8] , \Term[3][7] , 
        \Term[3][6] , \Term[3][5] , \Term[3][4] , \Term[3][3] , \Term[3][2] , 
        \Term[3][1] , \Term[3][0] }) );
  MUX_SHIFT_NB16_N_sh8 mux_map_4 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel(B[9:7]), .AS(OP[4]), .B({
        \Term[4][31] , \Term[4][30] , \Term[4][29] , \Term[4][28] , 
        \Term[4][27] , \Term[4][26] , \Term[4][25] , \Term[4][24] , 
        \Term[4][23] , \Term[4][22] , \Term[4][21] , \Term[4][20] , 
        \Term[4][19] , \Term[4][18] , \Term[4][17] , \Term[4][16] , 
        \Term[4][15] , \Term[4][14] , \Term[4][13] , \Term[4][12] , 
        \Term[4][11] , \Term[4][10] , \Term[4][9] , \Term[4][8] , \Term[4][7] , 
        \Term[4][6] , \Term[4][5] , \Term[4][4] , \Term[4][3] , \Term[4][2] , 
        \Term[4][1] , \Term[4][0] }) );
  MUX_SHIFT_NB16_N_sh10 mux_map_5 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel(B[11:9]), .AS(OP[5]), .B({
        \Term[5][31] , \Term[5][30] , \Term[5][29] , \Term[5][28] , 
        \Term[5][27] , \Term[5][26] , \Term[5][25] , \Term[5][24] , 
        \Term[5][23] , \Term[5][22] , \Term[5][21] , \Term[5][20] , 
        \Term[5][19] , \Term[5][18] , \Term[5][17] , \Term[5][16] , 
        \Term[5][15] , \Term[5][14] , \Term[5][13] , \Term[5][12] , 
        \Term[5][11] , \Term[5][10] , \Term[5][9] , \Term[5][8] , \Term[5][7] , 
        \Term[5][6] , \Term[5][5] , \Term[5][4] , \Term[5][3] , \Term[5][2] , 
        \Term[5][1] , \Term[5][0] }) );
  MUX_SHIFT_NB16_N_sh12 mux_map_6 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel(B[13:11]), .AS(OP[6]), .B({
        \Term[6][31] , \Term[6][30] , \Term[6][29] , \Term[6][28] , 
        \Term[6][27] , \Term[6][26] , \Term[6][25] , \Term[6][24] , 
        \Term[6][23] , \Term[6][22] , \Term[6][21] , \Term[6][20] , 
        \Term[6][19] , \Term[6][18] , \Term[6][17] , \Term[6][16] , 
        \Term[6][15] , \Term[6][14] , \Term[6][13] , \Term[6][12] , 
        \Term[6][11] , \Term[6][10] , \Term[6][9] , \Term[6][8] , \Term[6][7] , 
        \Term[6][6] , \Term[6][5] , \Term[6][4] , \Term[6][3] , \Term[6][2] , 
        \Term[6][1] , \Term[6][0] }) );
  MUX_SHIFT_NB16_N_sh14 mux_map_7 ( .A({n16, n15, n14, n13, n12, n11, n10, n9, 
        n8, n7, n6, n5, n4, n3, n2, n1}), .sel(B[15:13]), .AS(OP[7]), .B({
        \Term[7][31] , \Term[7][30] , \Term[7][29] , \Term[7][28] , 
        \Term[7][27] , \Term[7][26] , \Term[7][25] , \Term[7][24] , 
        \Term[7][23] , \Term[7][22] , \Term[7][21] , \Term[7][20] , 
        \Term[7][19] , \Term[7][18] , \Term[7][17] , \Term[7][16] , 
        \Term[7][15] , \Term[7][14] , \Term[7][13] , \Term[7][12] , 
        \Term[7][11] , \Term[7][10] , \Term[7][9] , \Term[7][8] , \Term[7][7] , 
        \Term[7][6] , \Term[7][5] , \Term[7][4] , \Term[7][3] , \Term[7][2] , 
        \Term[7][1] , \Term[7][0] }) );
  p4addgen_NB32_CW4_8 adder_0 ( .A({\Term[0][31] , \Term[0][30] , 
        \Term[0][29] , \Term[0][28] , \Term[0][27] , \Term[0][26] , 
        \Term[0][25] , \Term[0][24] , \Term[0][23] , \Term[0][22] , 
        \Term[0][21] , \Term[0][20] , \Term[0][19] , \Term[0][18] , 
        \Term[0][17] , \Term[0][16] , \Term[0][15] , \Term[0][14] , 
        \Term[0][13] , \Term[0][12] , \Term[0][11] , \Term[0][10] , 
        \Term[0][9] , \Term[0][8] , \Term[0][7] , \Term[0][6] , \Term[0][5] , 
        \Term[0][4] , \Term[0][3] , \Term[0][2] , \Term[0][1] , \Term[0][0] }), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Ci(OP[0]), 
        .S({\Res[0][31] , \Res[0][30] , \Res[0][29] , \Res[0][28] , 
        \Res[0][27] , \Res[0][26] , \Res[0][25] , \Res[0][24] , \Res[0][23] , 
        \Res[0][22] , \Res[0][21] , \Res[0][20] , \Res[0][19] , \Res[0][18] , 
        \Res[0][17] , \Res[0][16] , \Res[0][15] , \Res[0][14] , \Res[0][13] , 
        \Res[0][12] , \Res[0][11] , \Res[0][10] , \Res[0][9] , \Res[0][8] , 
        \Res[0][7] , \Res[0][6] , \Res[0][5] , \Res[0][4] , \Res[0][3] , 
        \Res[0][2] , \Res[0][1] , \Res[0][0] }) );
  p4addgen_NB32_CW4_7 add_map_1 ( .A({\Term[1][31] , \Term[1][30] , 
        \Term[1][29] , \Term[1][28] , \Term[1][27] , \Term[1][26] , 
        \Term[1][25] , \Term[1][24] , \Term[1][23] , \Term[1][22] , 
        \Term[1][21] , \Term[1][20] , \Term[1][19] , \Term[1][18] , 
        \Term[1][17] , \Term[1][16] , \Term[1][15] , \Term[1][14] , 
        \Term[1][13] , \Term[1][12] , \Term[1][11] , \Term[1][10] , 
        \Term[1][9] , \Term[1][8] , \Term[1][7] , \Term[1][6] , \Term[1][5] , 
        \Term[1][4] , \Term[1][3] , \Term[1][2] , \Term[1][1] , \Term[1][0] }), 
        .B({\Res[0][31] , \Res[0][30] , \Res[0][29] , \Res[0][28] , 
        \Res[0][27] , \Res[0][26] , \Res[0][25] , \Res[0][24] , \Res[0][23] , 
        \Res[0][22] , \Res[0][21] , \Res[0][20] , \Res[0][19] , \Res[0][18] , 
        \Res[0][17] , \Res[0][16] , \Res[0][15] , \Res[0][14] , \Res[0][13] , 
        \Res[0][12] , \Res[0][11] , \Res[0][10] , \Res[0][9] , \Res[0][8] , 
        \Res[0][7] , \Res[0][6] , \Res[0][5] , \Res[0][4] , \Res[0][3] , 
        \Res[0][2] , \Res[0][1] , \Res[0][0] }), .Ci(OP[1]), .S({\Res[1][31] , 
        \Res[1][30] , \Res[1][29] , \Res[1][28] , \Res[1][27] , \Res[1][26] , 
        \Res[1][25] , \Res[1][24] , \Res[1][23] , \Res[1][22] , \Res[1][21] , 
        \Res[1][20] , \Res[1][19] , \Res[1][18] , \Res[1][17] , \Res[1][16] , 
        \Res[1][15] , \Res[1][14] , \Res[1][13] , \Res[1][12] , \Res[1][11] , 
        \Res[1][10] , \Res[1][9] , \Res[1][8] , \Res[1][7] , \Res[1][6] , 
        \Res[1][5] , \Res[1][4] , \Res[1][3] , \Res[1][2] , \Res[1][1] , 
        \Res[1][0] }) );
  p4addgen_NB32_CW4_6 add_map_2 ( .A({\Term[2][31] , \Term[2][30] , 
        \Term[2][29] , \Term[2][28] , \Term[2][27] , \Term[2][26] , 
        \Term[2][25] , \Term[2][24] , \Term[2][23] , \Term[2][22] , 
        \Term[2][21] , \Term[2][20] , \Term[2][19] , \Term[2][18] , 
        \Term[2][17] , \Term[2][16] , \Term[2][15] , \Term[2][14] , 
        \Term[2][13] , \Term[2][12] , \Term[2][11] , \Term[2][10] , 
        \Term[2][9] , \Term[2][8] , \Term[2][7] , \Term[2][6] , \Term[2][5] , 
        \Term[2][4] , \Term[2][3] , \Term[2][2] , \Term[2][1] , \Term[2][0] }), 
        .B({\Res[1][31] , \Res[1][30] , \Res[1][29] , \Res[1][28] , 
        \Res[1][27] , \Res[1][26] , \Res[1][25] , \Res[1][24] , \Res[1][23] , 
        \Res[1][22] , \Res[1][21] , \Res[1][20] , \Res[1][19] , \Res[1][18] , 
        \Res[1][17] , \Res[1][16] , \Res[1][15] , \Res[1][14] , \Res[1][13] , 
        \Res[1][12] , \Res[1][11] , \Res[1][10] , \Res[1][9] , \Res[1][8] , 
        \Res[1][7] , \Res[1][6] , \Res[1][5] , \Res[1][4] , \Res[1][3] , 
        \Res[1][2] , \Res[1][1] , \Res[1][0] }), .Ci(OP[2]), .S({\Res[2][31] , 
        \Res[2][30] , \Res[2][29] , \Res[2][28] , \Res[2][27] , \Res[2][26] , 
        \Res[2][25] , \Res[2][24] , \Res[2][23] , \Res[2][22] , \Res[2][21] , 
        \Res[2][20] , \Res[2][19] , \Res[2][18] , \Res[2][17] , \Res[2][16] , 
        \Res[2][15] , \Res[2][14] , \Res[2][13] , \Res[2][12] , \Res[2][11] , 
        \Res[2][10] , \Res[2][9] , \Res[2][8] , \Res[2][7] , \Res[2][6] , 
        \Res[2][5] , \Res[2][4] , \Res[2][3] , \Res[2][2] , \Res[2][1] , 
        \Res[2][0] }) );
  p4addgen_NB32_CW4_5 add_map_3 ( .A({\Term[3][31] , \Term[3][30] , 
        \Term[3][29] , \Term[3][28] , \Term[3][27] , \Term[3][26] , 
        \Term[3][25] , \Term[3][24] , \Term[3][23] , \Term[3][22] , 
        \Term[3][21] , \Term[3][20] , \Term[3][19] , \Term[3][18] , 
        \Term[3][17] , \Term[3][16] , \Term[3][15] , \Term[3][14] , 
        \Term[3][13] , \Term[3][12] , \Term[3][11] , \Term[3][10] , 
        \Term[3][9] , \Term[3][8] , \Term[3][7] , \Term[3][6] , \Term[3][5] , 
        \Term[3][4] , \Term[3][3] , \Term[3][2] , \Term[3][1] , \Term[3][0] }), 
        .B({\Res[2][31] , \Res[2][30] , \Res[2][29] , \Res[2][28] , 
        \Res[2][27] , \Res[2][26] , \Res[2][25] , \Res[2][24] , \Res[2][23] , 
        \Res[2][22] , \Res[2][21] , \Res[2][20] , \Res[2][19] , \Res[2][18] , 
        \Res[2][17] , \Res[2][16] , \Res[2][15] , \Res[2][14] , \Res[2][13] , 
        \Res[2][12] , \Res[2][11] , \Res[2][10] , \Res[2][9] , \Res[2][8] , 
        \Res[2][7] , \Res[2][6] , \Res[2][5] , \Res[2][4] , \Res[2][3] , 
        \Res[2][2] , \Res[2][1] , \Res[2][0] }), .Ci(OP[3]), .S({\Res[3][31] , 
        \Res[3][30] , \Res[3][29] , \Res[3][28] , \Res[3][27] , \Res[3][26] , 
        \Res[3][25] , \Res[3][24] , \Res[3][23] , \Res[3][22] , \Res[3][21] , 
        \Res[3][20] , \Res[3][19] , \Res[3][18] , \Res[3][17] , \Res[3][16] , 
        \Res[3][15] , \Res[3][14] , \Res[3][13] , \Res[3][12] , \Res[3][11] , 
        \Res[3][10] , \Res[3][9] , \Res[3][8] , \Res[3][7] , \Res[3][6] , 
        \Res[3][5] , \Res[3][4] , \Res[3][3] , \Res[3][2] , \Res[3][1] , 
        \Res[3][0] }) );
  p4addgen_NB32_CW4_4 add_map_4 ( .A({\Term[4][31] , \Term[4][30] , 
        \Term[4][29] , \Term[4][28] , \Term[4][27] , \Term[4][26] , 
        \Term[4][25] , \Term[4][24] , \Term[4][23] , \Term[4][22] , 
        \Term[4][21] , \Term[4][20] , \Term[4][19] , \Term[4][18] , 
        \Term[4][17] , \Term[4][16] , \Term[4][15] , \Term[4][14] , 
        \Term[4][13] , \Term[4][12] , \Term[4][11] , \Term[4][10] , 
        \Term[4][9] , \Term[4][8] , \Term[4][7] , \Term[4][6] , \Term[4][5] , 
        \Term[4][4] , \Term[4][3] , \Term[4][2] , \Term[4][1] , \Term[4][0] }), 
        .B({\Res[3][31] , \Res[3][30] , \Res[3][29] , \Res[3][28] , 
        \Res[3][27] , \Res[3][26] , \Res[3][25] , \Res[3][24] , \Res[3][23] , 
        \Res[3][22] , \Res[3][21] , \Res[3][20] , \Res[3][19] , \Res[3][18] , 
        \Res[3][17] , \Res[3][16] , \Res[3][15] , \Res[3][14] , \Res[3][13] , 
        \Res[3][12] , \Res[3][11] , \Res[3][10] , \Res[3][9] , \Res[3][8] , 
        \Res[3][7] , \Res[3][6] , \Res[3][5] , \Res[3][4] , \Res[3][3] , 
        \Res[3][2] , \Res[3][1] , \Res[3][0] }), .Ci(OP[4]), .S({\Res[4][31] , 
        \Res[4][30] , \Res[4][29] , \Res[4][28] , \Res[4][27] , \Res[4][26] , 
        \Res[4][25] , \Res[4][24] , \Res[4][23] , \Res[4][22] , \Res[4][21] , 
        \Res[4][20] , \Res[4][19] , \Res[4][18] , \Res[4][17] , \Res[4][16] , 
        \Res[4][15] , \Res[4][14] , \Res[4][13] , \Res[4][12] , \Res[4][11] , 
        \Res[4][10] , \Res[4][9] , \Res[4][8] , \Res[4][7] , \Res[4][6] , 
        \Res[4][5] , \Res[4][4] , \Res[4][3] , \Res[4][2] , \Res[4][1] , 
        \Res[4][0] }) );
  p4addgen_NB32_CW4_3 add_map_5 ( .A({\Term[5][31] , \Term[5][30] , 
        \Term[5][29] , \Term[5][28] , \Term[5][27] , \Term[5][26] , 
        \Term[5][25] , \Term[5][24] , \Term[5][23] , \Term[5][22] , 
        \Term[5][21] , \Term[5][20] , \Term[5][19] , \Term[5][18] , 
        \Term[5][17] , \Term[5][16] , \Term[5][15] , \Term[5][14] , 
        \Term[5][13] , \Term[5][12] , \Term[5][11] , \Term[5][10] , 
        \Term[5][9] , \Term[5][8] , \Term[5][7] , \Term[5][6] , \Term[5][5] , 
        \Term[5][4] , \Term[5][3] , \Term[5][2] , \Term[5][1] , \Term[5][0] }), 
        .B({\Res[4][31] , \Res[4][30] , \Res[4][29] , \Res[4][28] , 
        \Res[4][27] , \Res[4][26] , \Res[4][25] , \Res[4][24] , \Res[4][23] , 
        \Res[4][22] , \Res[4][21] , \Res[4][20] , \Res[4][19] , \Res[4][18] , 
        \Res[4][17] , \Res[4][16] , \Res[4][15] , \Res[4][14] , \Res[4][13] , 
        \Res[4][12] , \Res[4][11] , \Res[4][10] , \Res[4][9] , \Res[4][8] , 
        \Res[4][7] , \Res[4][6] , \Res[4][5] , \Res[4][4] , \Res[4][3] , 
        \Res[4][2] , \Res[4][1] , \Res[4][0] }), .Ci(OP[5]), .S({\Res[5][31] , 
        \Res[5][30] , \Res[5][29] , \Res[5][28] , \Res[5][27] , \Res[5][26] , 
        \Res[5][25] , \Res[5][24] , \Res[5][23] , \Res[5][22] , \Res[5][21] , 
        \Res[5][20] , \Res[5][19] , \Res[5][18] , \Res[5][17] , \Res[5][16] , 
        \Res[5][15] , \Res[5][14] , \Res[5][13] , \Res[5][12] , \Res[5][11] , 
        \Res[5][10] , \Res[5][9] , \Res[5][8] , \Res[5][7] , \Res[5][6] , 
        \Res[5][5] , \Res[5][4] , \Res[5][3] , \Res[5][2] , \Res[5][1] , 
        \Res[5][0] }) );
  p4addgen_NB32_CW4_2 add_map_6 ( .A({\Term[6][31] , \Term[6][30] , 
        \Term[6][29] , \Term[6][28] , \Term[6][27] , \Term[6][26] , 
        \Term[6][25] , \Term[6][24] , \Term[6][23] , \Term[6][22] , 
        \Term[6][21] , \Term[6][20] , \Term[6][19] , \Term[6][18] , 
        \Term[6][17] , \Term[6][16] , \Term[6][15] , \Term[6][14] , 
        \Term[6][13] , \Term[6][12] , \Term[6][11] , \Term[6][10] , 
        \Term[6][9] , \Term[6][8] , \Term[6][7] , \Term[6][6] , \Term[6][5] , 
        \Term[6][4] , \Term[6][3] , \Term[6][2] , \Term[6][1] , \Term[6][0] }), 
        .B({\Res[5][31] , \Res[5][30] , \Res[5][29] , \Res[5][28] , 
        \Res[5][27] , \Res[5][26] , \Res[5][25] , \Res[5][24] , \Res[5][23] , 
        \Res[5][22] , \Res[5][21] , \Res[5][20] , \Res[5][19] , \Res[5][18] , 
        \Res[5][17] , \Res[5][16] , \Res[5][15] , \Res[5][14] , \Res[5][13] , 
        \Res[5][12] , \Res[5][11] , \Res[5][10] , \Res[5][9] , \Res[5][8] , 
        \Res[5][7] , \Res[5][6] , \Res[5][5] , \Res[5][4] , \Res[5][3] , 
        \Res[5][2] , \Res[5][1] , \Res[5][0] }), .Ci(OP[6]), .S({\Res[6][31] , 
        \Res[6][30] , \Res[6][29] , \Res[6][28] , \Res[6][27] , \Res[6][26] , 
        \Res[6][25] , \Res[6][24] , \Res[6][23] , \Res[6][22] , \Res[6][21] , 
        \Res[6][20] , \Res[6][19] , \Res[6][18] , \Res[6][17] , \Res[6][16] , 
        \Res[6][15] , \Res[6][14] , \Res[6][13] , \Res[6][12] , \Res[6][11] , 
        \Res[6][10] , \Res[6][9] , \Res[6][8] , \Res[6][7] , \Res[6][6] , 
        \Res[6][5] , \Res[6][4] , \Res[6][3] , \Res[6][2] , \Res[6][1] , 
        \Res[6][0] }) );
  p4addgen_NB32_CW4_1 add_map_7 ( .A({\Term[7][31] , \Term[7][30] , 
        \Term[7][29] , \Term[7][28] , \Term[7][27] , \Term[7][26] , 
        \Term[7][25] , \Term[7][24] , \Term[7][23] , \Term[7][22] , 
        \Term[7][21] , \Term[7][20] , \Term[7][19] , \Term[7][18] , 
        \Term[7][17] , \Term[7][16] , \Term[7][15] , \Term[7][14] , 
        \Term[7][13] , \Term[7][12] , \Term[7][11] , \Term[7][10] , 
        \Term[7][9] , \Term[7][8] , \Term[7][7] , \Term[7][6] , \Term[7][5] , 
        \Term[7][4] , \Term[7][3] , \Term[7][2] , \Term[7][1] , \Term[7][0] }), 
        .B({\Res[6][31] , \Res[6][30] , \Res[6][29] , \Res[6][28] , 
        \Res[6][27] , \Res[6][26] , \Res[6][25] , \Res[6][24] , \Res[6][23] , 
        \Res[6][22] , \Res[6][21] , \Res[6][20] , \Res[6][19] , \Res[6][18] , 
        \Res[6][17] , \Res[6][16] , \Res[6][15] , \Res[6][14] , \Res[6][13] , 
        \Res[6][12] , \Res[6][11] , \Res[6][10] , \Res[6][9] , \Res[6][8] , 
        \Res[6][7] , \Res[6][6] , \Res[6][5] , \Res[6][4] , \Res[6][3] , 
        \Res[6][2] , \Res[6][1] , \Res[6][0] }), .Ci(OP[7]), .S(C) );
  BUF_X1 U2 ( .A(A[15]), .Z(n16) );
endmodule


module p4addgen_NB32_CW4_0 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] carry_sh;

  CSTgen_CW4_NB32_0 sparse_tree ( .A(A), .B(B), .Ci(Ci), .C({Co, carry_sh}) );
  sum_gen_Nrca4_NB32_0 carry_sel ( .A(A), .B(B), .Ci({carry_sh, Ci}), .S(S) );
endmodule


module MUX31_generic_NB32_1 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n153, n154, n155, n157, n158, n159,
         n160, n161, n162, n163, n164, n165;

  INV_X2 U8 ( .A(n40), .ZN(Y[6]) );
  INV_X2 U54 ( .A(n63), .ZN(Y[14]) );
  INV_X2 U58 ( .A(n65), .ZN(Y[12]) );
  INV_X1 U2 ( .A(n57), .ZN(Y[1]) );
  OR3_X2 U3 ( .A1(n153), .A2(n154), .A3(n155), .ZN(Y[9]) );
  AND2_X1 U4 ( .A1(C[9]), .A2(n165), .ZN(n153) );
  AND2_X1 U5 ( .A1(B[9]), .A2(n162), .ZN(n154) );
  AND2_X1 U6 ( .A1(A[9]), .A2(n159), .ZN(n155) );
  BUF_X2 U7 ( .A(n35), .Z(n163) );
  BUF_X2 U9 ( .A(n36), .Z(n161) );
  BUF_X2 U10 ( .A(n35), .Z(n164) );
  BUF_X1 U11 ( .A(n37), .Z(n159) );
  BUF_X2 U12 ( .A(n37), .Z(n158) );
  INV_X1 U13 ( .A(SEL[0]), .ZN(n69) );
  INV_X1 U14 ( .A(n44), .ZN(Y[31]) );
  INV_X1 U15 ( .A(n42), .ZN(Y[4]) );
  INV_X1 U16 ( .A(n46), .ZN(Y[2]) );
  INV_X1 U17 ( .A(n43), .ZN(Y[3]) );
  INV_X1 U18 ( .A(n39), .ZN(Y[7]) );
  INV_X1 U19 ( .A(n38), .ZN(Y[8]) );
  INV_X1 U20 ( .A(n66), .ZN(Y[11]) );
  INV_X1 U21 ( .A(n64), .ZN(Y[13]) );
  INV_X1 U22 ( .A(n62), .ZN(Y[15]) );
  INV_X1 U23 ( .A(n59), .ZN(Y[18]) );
  INV_X1 U24 ( .A(n61), .ZN(Y[16]) );
  INV_X1 U25 ( .A(n60), .ZN(Y[17]) );
  INV_X1 U26 ( .A(n58), .ZN(Y[19]) );
  INV_X1 U27 ( .A(n54), .ZN(Y[22]) );
  INV_X1 U28 ( .A(n52), .ZN(Y[24]) );
  INV_X1 U29 ( .A(n56), .ZN(Y[20]) );
  INV_X1 U30 ( .A(n51), .ZN(Y[25]) );
  INV_X1 U31 ( .A(n53), .ZN(Y[23]) );
  INV_X1 U32 ( .A(n47), .ZN(Y[29]) );
  INV_X1 U33 ( .A(n48), .ZN(Y[28]) );
  AOI222_X1 U34 ( .A1(C[28]), .A2(n164), .B1(B[28]), .B2(n161), .C1(A[28]), 
        .C2(n157), .ZN(n48) );
  INV_X1 U35 ( .A(n50), .ZN(Y[26]) );
  AOI222_X1 U36 ( .A1(C[26]), .A2(n164), .B1(B[26]), .B2(n161), .C1(A[26]), 
        .C2(n157), .ZN(n50) );
  INV_X1 U37 ( .A(n55), .ZN(Y[21]) );
  AOI222_X1 U38 ( .A1(C[21]), .A2(n164), .B1(B[21]), .B2(n161), .C1(A[21]), 
        .C2(n157), .ZN(n55) );
  INV_X1 U39 ( .A(n49), .ZN(Y[27]) );
  AOI222_X1 U40 ( .A1(C[27]), .A2(n164), .B1(B[27]), .B2(n161), .C1(A[27]), 
        .C2(n157), .ZN(n49) );
  INV_X1 U41 ( .A(n45), .ZN(Y[30]) );
  AOI222_X1 U42 ( .A1(C[30]), .A2(n164), .B1(B[30]), .B2(n161), .C1(A[30]), 
        .C2(n157), .ZN(n45) );
  AOI222_X1 U43 ( .A1(C[29]), .A2(n164), .B1(B[29]), .B2(n161), .C1(A[29]), 
        .C2(n158), .ZN(n47) );
  AOI222_X1 U44 ( .A1(C[24]), .A2(n164), .B1(B[24]), .B2(n161), .C1(A[24]), 
        .C2(n158), .ZN(n52) );
  AOI222_X1 U45 ( .A1(C[25]), .A2(n164), .B1(B[25]), .B2(n161), .C1(A[25]), 
        .C2(n158), .ZN(n51) );
  AOI222_X1 U46 ( .A1(C[20]), .A2(n164), .B1(B[20]), .B2(n161), .C1(A[20]), 
        .C2(n158), .ZN(n56) );
  AOI222_X1 U47 ( .A1(C[22]), .A2(n164), .B1(B[22]), .B2(n161), .C1(A[22]), 
        .C2(n158), .ZN(n54) );
  AOI222_X1 U48 ( .A1(C[23]), .A2(n164), .B1(B[23]), .B2(n161), .C1(A[23]), 
        .C2(n158), .ZN(n53) );
  AOI222_X1 U49 ( .A1(C[2]), .A2(n164), .B1(B[2]), .B2(n161), .C1(A[2]), .C2(
        n158), .ZN(n46) );
  AOI222_X1 U50 ( .A1(C[14]), .A2(n163), .B1(B[14]), .B2(n160), .C1(A[14]), 
        .C2(n158), .ZN(n63) );
  INV_X1 U51 ( .A(n41), .ZN(Y[5]) );
  INV_X1 U52 ( .A(n67), .ZN(Y[10]) );
  BUF_X2 U53 ( .A(n36), .Z(n160) );
  BUF_X2 U55 ( .A(n35), .Z(n165) );
  AOI222_X1 U56 ( .A1(C[31]), .A2(n165), .B1(B[31]), .B2(n162), .C1(A[31]), 
        .C2(n157), .ZN(n44) );
  AOI222_X1 U57 ( .A1(C[8]), .A2(n165), .B1(B[8]), .B2(n162), .C1(A[8]), .C2(
        n157), .ZN(n38) );
  AOI222_X1 U59 ( .A1(C[4]), .A2(n165), .B1(B[4]), .B2(n162), .C1(A[4]), .C2(
        n158), .ZN(n42) );
  AOI222_X1 U60 ( .A1(C[5]), .A2(n165), .B1(B[5]), .B2(n162), .C1(A[5]), .C2(
        n158), .ZN(n41) );
  AOI222_X1 U61 ( .A1(C[3]), .A2(n165), .B1(B[3]), .B2(n162), .C1(A[3]), .C2(
        n159), .ZN(n43) );
  AOI222_X1 U62 ( .A1(C[7]), .A2(n165), .B1(B[7]), .B2(n162), .C1(A[7]), .C2(
        n159), .ZN(n39) );
  BUF_X2 U63 ( .A(n36), .Z(n162) );
  AOI222_X1 U64 ( .A1(C[6]), .A2(n165), .B1(B[6]), .B2(n162), .C1(A[6]), .C2(
        n159), .ZN(n40) );
  AOI222_X1 U65 ( .A1(C[16]), .A2(n163), .B1(B[16]), .B2(n160), .C1(A[16]), 
        .C2(n157), .ZN(n61) );
  AOI222_X1 U66 ( .A1(C[18]), .A2(n163), .B1(B[18]), .B2(n160), .C1(A[18]), 
        .C2(n157), .ZN(n59) );
  AOI222_X1 U67 ( .A1(C[11]), .A2(n163), .B1(B[11]), .B2(n160), .C1(A[11]), 
        .C2(n157), .ZN(n66) );
  AOI222_X1 U68 ( .A1(C[17]), .A2(n163), .B1(B[17]), .B2(n160), .C1(A[17]), 
        .C2(n157), .ZN(n60) );
  AOI222_X1 U69 ( .A1(C[19]), .A2(n163), .B1(B[19]), .B2(n160), .C1(A[19]), 
        .C2(n157), .ZN(n58) );
  AOI222_X1 U70 ( .A1(C[15]), .A2(n163), .B1(B[15]), .B2(n160), .C1(A[15]), 
        .C2(n158), .ZN(n62) );
  AOI222_X1 U71 ( .A1(C[13]), .A2(n163), .B1(B[13]), .B2(n160), .C1(A[13]), 
        .C2(n157), .ZN(n64) );
  AOI222_X1 U72 ( .A1(C[10]), .A2(n163), .B1(B[10]), .B2(n160), .C1(A[10]), 
        .C2(n159), .ZN(n67) );
  AOI222_X1 U73 ( .A1(C[12]), .A2(n163), .B1(B[12]), .B2(n160), .C1(A[12]), 
        .C2(n158), .ZN(n65) );
  AOI222_X1 U74 ( .A1(C[1]), .A2(n163), .B1(B[1]), .B2(n160), .C1(A[1]), .C2(
        n159), .ZN(n57) );
  AOI222_X1 U75 ( .A1(C[0]), .A2(n163), .B1(B[0]), .B2(n160), .C1(A[0]), .C2(
        n159), .ZN(n68) );
  BUF_X2 U76 ( .A(n37), .Z(n157) );
  INV_X1 U77 ( .A(n68), .ZN(Y[0]) );
  AND2_X1 U78 ( .A1(SEL[1]), .A2(n69), .ZN(n35) );
  NOR2_X1 U79 ( .A1(n69), .A2(SEL[1]), .ZN(n36) );
  NOR2_X1 U80 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n37) );
endmodule


module MUX31_generic_NB32_0 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n159, n160, n161, n162, n163,
         n164, n165, n166, n167;

  BUF_X2 U2 ( .A(n35), .Z(n165) );
  INV_X1 U3 ( .A(SEL[0]), .ZN(n69) );
  BUF_X2 U4 ( .A(n36), .Z(n164) );
  BUF_X2 U5 ( .A(n36), .Z(n163) );
  BUF_X2 U6 ( .A(n37), .Z(n160) );
  CLKBUF_X3 U7 ( .A(n35), .Z(n166) );
  BUF_X2 U8 ( .A(n35), .Z(n167) );
  BUF_X1 U9 ( .A(n36), .Z(n162) );
  BUF_X1 U10 ( .A(n37), .Z(n159) );
  INV_X1 U11 ( .A(n65), .ZN(Y[12]) );
  INV_X1 U12 ( .A(n42), .ZN(Y[4]) );
  INV_X1 U13 ( .A(n63), .ZN(Y[14]) );
  INV_X1 U14 ( .A(n44), .ZN(Y[31]) );
  AOI222_X1 U15 ( .A1(C[31]), .A2(n167), .B1(B[31]), .B2(n164), .C1(A[31]), 
        .C2(n161), .ZN(n44) );
  INV_X1 U16 ( .A(n40), .ZN(Y[6]) );
  INV_X1 U17 ( .A(n60), .ZN(Y[17]) );
  INV_X1 U18 ( .A(n59), .ZN(Y[18]) );
  INV_X1 U19 ( .A(n61), .ZN(Y[16]) );
  INV_X1 U20 ( .A(n50), .ZN(Y[26]) );
  INV_X1 U21 ( .A(n54), .ZN(Y[22]) );
  INV_X1 U22 ( .A(n67), .ZN(Y[10]) );
  INV_X1 U23 ( .A(n45), .ZN(Y[30]) );
  INV_X1 U24 ( .A(n51), .ZN(Y[25]) );
  AOI222_X1 U25 ( .A1(C[25]), .A2(n166), .B1(B[25]), .B2(n164), .C1(A[25]), 
        .C2(n161), .ZN(n51) );
  INV_X1 U26 ( .A(n48), .ZN(Y[28]) );
  AOI222_X1 U27 ( .A1(C[28]), .A2(n166), .B1(B[28]), .B2(n164), .C1(A[28]), 
        .C2(n161), .ZN(n48) );
  INV_X1 U28 ( .A(n55), .ZN(Y[21]) );
  AOI222_X1 U29 ( .A1(C[21]), .A2(n166), .B1(B[21]), .B2(n163), .C1(A[21]), 
        .C2(n161), .ZN(n55) );
  INV_X1 U30 ( .A(n52), .ZN(Y[24]) );
  AOI222_X1 U31 ( .A1(C[24]), .A2(n166), .B1(B[24]), .B2(n164), .C1(A[24]), 
        .C2(n161), .ZN(n52) );
  INV_X1 U32 ( .A(n49), .ZN(Y[27]) );
  INV_X1 U33 ( .A(n53), .ZN(Y[23]) );
  INV_X1 U34 ( .A(n47), .ZN(Y[29]) );
  INV_X1 U35 ( .A(n56), .ZN(Y[20]) );
  AOI222_X1 U36 ( .A1(C[20]), .A2(n166), .B1(B[20]), .B2(n164), .C1(A[20]), 
        .C2(n161), .ZN(n56) );
  INV_X1 U37 ( .A(n58), .ZN(Y[19]) );
  INV_X1 U38 ( .A(n62), .ZN(Y[15]) );
  AOI222_X1 U39 ( .A1(C[8]), .A2(n167), .B1(B[8]), .B2(n164), .C1(A[8]), .C2(
        n161), .ZN(n38) );
  BUF_X2 U40 ( .A(n37), .Z(n161) );
  INV_X1 U41 ( .A(n38), .ZN(Y[8]) );
  AOI222_X1 U42 ( .A1(C[4]), .A2(n167), .B1(B[4]), .B2(n162), .C1(A[4]), .C2(
        n159), .ZN(n42) );
  AOI222_X1 U43 ( .A1(C[3]), .A2(n167), .B1(B[3]), .B2(n162), .C1(A[3]), .C2(
        n159), .ZN(n43) );
  AOI222_X1 U44 ( .A1(C[6]), .A2(n167), .B1(B[6]), .B2(n162), .C1(A[6]), .C2(
        n159), .ZN(n40) );
  AOI222_X1 U45 ( .A1(C[30]), .A2(n166), .B1(B[30]), .B2(n163), .C1(A[30]), 
        .C2(n160), .ZN(n45) );
  AOI222_X1 U46 ( .A1(C[29]), .A2(n166), .B1(B[29]), .B2(n163), .C1(A[29]), 
        .C2(n160), .ZN(n47) );
  AOI222_X1 U47 ( .A1(C[26]), .A2(n166), .B1(B[26]), .B2(n163), .C1(A[26]), 
        .C2(n160), .ZN(n50) );
  AOI222_X1 U48 ( .A1(C[27]), .A2(n166), .B1(B[27]), .B2(n163), .C1(A[27]), 
        .C2(n160), .ZN(n49) );
  AOI222_X1 U49 ( .A1(C[22]), .A2(n166), .B1(B[22]), .B2(n163), .C1(A[22]), 
        .C2(n160), .ZN(n54) );
  AOI222_X1 U50 ( .A1(C[23]), .A2(n166), .B1(B[23]), .B2(n164), .C1(A[23]), 
        .C2(n160), .ZN(n53) );
  AOI222_X1 U51 ( .A1(C[2]), .A2(n166), .B1(B[2]), .B2(n162), .C1(A[2]), .C2(
        n160), .ZN(n46) );
  AOI222_X1 U52 ( .A1(C[5]), .A2(n167), .B1(B[5]), .B2(n164), .C1(A[5]), .C2(
        n160), .ZN(n41) );
  AOI222_X1 U53 ( .A1(C[9]), .A2(n167), .B1(B[9]), .B2(n164), .C1(A[9]), .C2(
        n160), .ZN(n34) );
  INV_X1 U54 ( .A(n34), .ZN(Y[9]) );
  INV_X1 U55 ( .A(n57), .ZN(Y[1]) );
  INV_X1 U56 ( .A(n46), .ZN(Y[2]) );
  INV_X1 U57 ( .A(n41), .ZN(Y[5]) );
  AOI222_X1 U58 ( .A1(C[16]), .A2(n165), .B1(B[16]), .B2(n163), .C1(A[16]), 
        .C2(n160), .ZN(n61) );
  AOI222_X1 U59 ( .A1(C[18]), .A2(n165), .B1(B[18]), .B2(n164), .C1(A[18]), 
        .C2(n161), .ZN(n59) );
  AOI222_X1 U60 ( .A1(C[15]), .A2(n165), .B1(B[15]), .B2(n163), .C1(A[15]), 
        .C2(n161), .ZN(n62) );
  AOI222_X1 U61 ( .A1(C[19]), .A2(n165), .B1(B[19]), .B2(n163), .C1(A[19]), 
        .C2(n161), .ZN(n58) );
  AOI222_X1 U62 ( .A1(C[17]), .A2(n165), .B1(B[17]), .B2(n163), .C1(A[17]), 
        .C2(n161), .ZN(n60) );
  AOI222_X1 U63 ( .A1(C[10]), .A2(n165), .B1(B[10]), .B2(n164), .C1(A[10]), 
        .C2(n161), .ZN(n67) );
  AOI222_X1 U64 ( .A1(C[13]), .A2(n165), .B1(B[13]), .B2(n163), .C1(A[13]), 
        .C2(n161), .ZN(n64) );
  AOI222_X1 U65 ( .A1(C[12]), .A2(n165), .B1(B[12]), .B2(n163), .C1(A[12]), 
        .C2(n159), .ZN(n65) );
  AOI222_X1 U66 ( .A1(C[14]), .A2(n165), .B1(B[14]), .B2(n162), .C1(A[14]), 
        .C2(n159), .ZN(n63) );
  AOI222_X1 U67 ( .A1(C[1]), .A2(n165), .B1(B[1]), .B2(n163), .C1(A[1]), .C2(
        n160), .ZN(n57) );
  AOI222_X1 U68 ( .A1(C[0]), .A2(n165), .B1(B[0]), .B2(n162), .C1(A[0]), .C2(
        n159), .ZN(n68) );
  AOI222_X1 U69 ( .A1(C[11]), .A2(n165), .B1(B[11]), .B2(n164), .C1(A[11]), 
        .C2(n160), .ZN(n66) );
  INV_X1 U70 ( .A(n66), .ZN(Y[11]) );
  INV_X1 U71 ( .A(n64), .ZN(Y[13]) );
  AOI222_X1 U72 ( .A1(C[7]), .A2(n167), .B1(B[7]), .B2(n163), .C1(A[7]), .C2(
        n161), .ZN(n39) );
  INV_X1 U73 ( .A(n39), .ZN(Y[7]) );
  INV_X1 U74 ( .A(n43), .ZN(Y[3]) );
  INV_X1 U75 ( .A(n68), .ZN(Y[0]) );
  AND2_X1 U76 ( .A1(SEL[1]), .A2(n69), .ZN(n35) );
  NOR2_X1 U77 ( .A1(n69), .A2(SEL[1]), .ZN(n36) );
  NOR2_X1 U78 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n37) );
endmodule


module MUX21_generic_NB32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77;

  INV_X1 U1 ( .A(n76), .ZN(n67) );
  BUF_X1 U2 ( .A(n77), .Z(n69) );
  BUF_X1 U3 ( .A(n77), .Z(n68) );
  BUF_X1 U4 ( .A(n74), .Z(n70) );
  BUF_X1 U5 ( .A(n68), .Z(n75) );
  BUF_X1 U6 ( .A(n73), .Z(n74) );
  BUF_X1 U7 ( .A(n77), .Z(n73) );
  BUF_X1 U8 ( .A(n77), .Z(n72) );
  BUF_X1 U9 ( .A(n77), .Z(n71) );
  BUF_X1 U10 ( .A(n77), .Z(n76) );
  INV_X1 U11 ( .A(SEL), .ZN(n77) );
  INV_X1 U12 ( .A(n63), .ZN(Y[12]) );
  AOI22_X1 U13 ( .A1(A[12]), .A2(n67), .B1(B[12]), .B2(n75), .ZN(n63) );
  INV_X1 U14 ( .A(n38), .ZN(Y[6]) );
  AOI22_X1 U15 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(n68), .ZN(n38) );
  INV_X1 U16 ( .A(n61), .ZN(Y[14]) );
  AOI22_X1 U17 ( .A1(A[14]), .A2(n67), .B1(B[14]), .B2(n74), .ZN(n61) );
  INV_X1 U18 ( .A(n42), .ZN(Y[31]) );
  AOI22_X1 U19 ( .A1(A[31]), .A2(SEL), .B1(B[31]), .B2(n69), .ZN(n42) );
  INV_X1 U20 ( .A(n40), .ZN(Y[4]) );
  AOI22_X1 U21 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(n69), .ZN(n40) );
  INV_X1 U22 ( .A(n39), .ZN(Y[5]) );
  AOI22_X1 U23 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(n69), .ZN(n39) );
  INV_X1 U24 ( .A(n44), .ZN(Y[2]) );
  AOI22_X1 U25 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n70), .ZN(n44) );
  INV_X1 U26 ( .A(n55), .ZN(Y[1]) );
  AOI22_X1 U27 ( .A1(A[1]), .A2(n67), .B1(B[1]), .B2(n73), .ZN(n55) );
  INV_X1 U28 ( .A(n41), .ZN(Y[3]) );
  AOI22_X1 U29 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(n69), .ZN(n41) );
  INV_X1 U30 ( .A(n37), .ZN(Y[7]) );
  AOI22_X1 U31 ( .A1(A[7]), .A2(n67), .B1(B[7]), .B2(n68), .ZN(n37) );
  INV_X1 U32 ( .A(n36), .ZN(Y[8]) );
  AOI22_X1 U33 ( .A1(A[8]), .A2(SEL), .B1(B[8]), .B2(n68), .ZN(n36) );
  INV_X1 U34 ( .A(n64), .ZN(Y[11]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n67), .B1(B[11]), .B2(n75), .ZN(n64) );
  INV_X1 U36 ( .A(n62), .ZN(Y[13]) );
  AOI22_X1 U37 ( .A1(A[13]), .A2(n67), .B1(B[13]), .B2(n74), .ZN(n62) );
  INV_X1 U38 ( .A(n65), .ZN(Y[10]) );
  AOI22_X1 U39 ( .A1(A[10]), .A2(n67), .B1(B[10]), .B2(n75), .ZN(n65) );
  INV_X1 U40 ( .A(n66), .ZN(Y[0]) );
  AOI22_X1 U41 ( .A1(A[0]), .A2(n67), .B1(B[0]), .B2(n75), .ZN(n66) );
  INV_X1 U42 ( .A(n60), .ZN(Y[15]) );
  AOI22_X1 U43 ( .A1(A[15]), .A2(n67), .B1(B[15]), .B2(n74), .ZN(n60) );
  AOI22_X1 U44 ( .A1(n67), .A2(A[9]), .B1(B[9]), .B2(n68), .ZN(n34) );
  INV_X1 U45 ( .A(n57), .ZN(Y[18]) );
  AOI22_X1 U46 ( .A1(A[18]), .A2(n67), .B1(B[18]), .B2(n73), .ZN(n57) );
  INV_X1 U47 ( .A(n59), .ZN(Y[16]) );
  AOI22_X1 U48 ( .A1(A[16]), .A2(n67), .B1(B[16]), .B2(n74), .ZN(n59) );
  INV_X1 U49 ( .A(n58), .ZN(Y[17]) );
  AOI22_X1 U50 ( .A1(A[17]), .A2(n67), .B1(B[17]), .B2(n73), .ZN(n58) );
  INV_X1 U51 ( .A(n56), .ZN(Y[19]) );
  AOI22_X1 U52 ( .A1(A[19]), .A2(n67), .B1(B[19]), .B2(n73), .ZN(n56) );
  INV_X1 U53 ( .A(n52), .ZN(Y[22]) );
  AOI22_X1 U54 ( .A1(A[22]), .A2(SEL), .B1(B[22]), .B2(n72), .ZN(n52) );
  INV_X1 U55 ( .A(n50), .ZN(Y[24]) );
  AOI22_X1 U56 ( .A1(A[24]), .A2(SEL), .B1(B[24]), .B2(n71), .ZN(n50) );
  INV_X1 U57 ( .A(n54), .ZN(Y[20]) );
  AOI22_X1 U58 ( .A1(A[20]), .A2(SEL), .B1(B[20]), .B2(n72), .ZN(n54) );
  INV_X1 U59 ( .A(n49), .ZN(Y[25]) );
  AOI22_X1 U60 ( .A1(A[25]), .A2(SEL), .B1(B[25]), .B2(n71), .ZN(n49) );
  INV_X1 U61 ( .A(n51), .ZN(Y[23]) );
  AOI22_X1 U62 ( .A1(A[23]), .A2(SEL), .B1(B[23]), .B2(n72), .ZN(n51) );
  INV_X1 U63 ( .A(n45), .ZN(Y[29]) );
  AOI22_X1 U64 ( .A1(A[29]), .A2(SEL), .B1(B[29]), .B2(n70), .ZN(n45) );
  INV_X1 U65 ( .A(n46), .ZN(Y[28]) );
  AOI22_X1 U66 ( .A1(A[28]), .A2(SEL), .B1(B[28]), .B2(n70), .ZN(n46) );
  INV_X1 U67 ( .A(n48), .ZN(Y[26]) );
  AOI22_X1 U68 ( .A1(A[26]), .A2(SEL), .B1(B[26]), .B2(n71), .ZN(n48) );
  INV_X1 U69 ( .A(n53), .ZN(Y[21]) );
  AOI22_X1 U70 ( .A1(A[21]), .A2(SEL), .B1(B[21]), .B2(n72), .ZN(n53) );
  INV_X1 U71 ( .A(n47), .ZN(Y[27]) );
  AOI22_X1 U72 ( .A1(A[27]), .A2(SEL), .B1(B[27]), .B2(n71), .ZN(n47) );
  INV_X1 U73 ( .A(n43), .ZN(Y[30]) );
  AOI22_X1 U74 ( .A1(A[30]), .A2(SEL), .B1(B[30]), .B2(n70), .ZN(n43) );
  INV_X1 U75 ( .A(n34), .ZN(Y[9]) );
endmodule


module MUX21_generic_NB32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75;

  BUF_X1 U1 ( .A(n75), .Z(n68) );
  BUF_X1 U2 ( .A(n75), .Z(n74) );
  BUF_X1 U3 ( .A(n75), .Z(n73) );
  BUF_X1 U4 ( .A(n72), .Z(n67) );
  BUF_X1 U5 ( .A(n74), .Z(n69) );
  BUF_X1 U6 ( .A(n75), .Z(n72) );
  BUF_X1 U7 ( .A(n75), .Z(n71) );
  BUF_X1 U8 ( .A(n75), .Z(n70) );
  INV_X1 U9 ( .A(SEL), .ZN(n75) );
  INV_X1 U10 ( .A(n63), .ZN(Y[12]) );
  INV_X1 U11 ( .A(n40), .ZN(Y[4]) );
  INV_X1 U12 ( .A(n61), .ZN(Y[14]) );
  INV_X1 U13 ( .A(n42), .ZN(Y[31]) );
  AOI22_X1 U14 ( .A1(A[31]), .A2(SEL), .B1(B[31]), .B2(n68), .ZN(n42) );
  INV_X1 U15 ( .A(n38), .ZN(Y[6]) );
  INV_X1 U16 ( .A(n44), .ZN(Y[2]) );
  INV_X1 U17 ( .A(n36), .ZN(Y[8]) );
  INV_X1 U18 ( .A(n58), .ZN(Y[17]) );
  AOI22_X1 U19 ( .A1(A[17]), .A2(SEL), .B1(B[17]), .B2(n72), .ZN(n58) );
  INV_X1 U20 ( .A(n64), .ZN(Y[11]) );
  INV_X1 U21 ( .A(n57), .ZN(Y[18]) );
  AOI22_X1 U22 ( .A1(A[18]), .A2(SEL), .B1(B[18]), .B2(n72), .ZN(n57) );
  INV_X1 U23 ( .A(n41), .ZN(Y[3]) );
  INV_X1 U24 ( .A(n59), .ZN(Y[16]) );
  AOI22_X1 U25 ( .A1(A[16]), .A2(SEL), .B1(B[16]), .B2(n73), .ZN(n59) );
  INV_X1 U26 ( .A(n48), .ZN(Y[26]) );
  AOI22_X1 U27 ( .A1(A[26]), .A2(SEL), .B1(B[26]), .B2(n70), .ZN(n48) );
  INV_X1 U28 ( .A(n52), .ZN(Y[22]) );
  AOI22_X1 U29 ( .A1(A[22]), .A2(SEL), .B1(B[22]), .B2(n71), .ZN(n52) );
  INV_X1 U30 ( .A(n55), .ZN(Y[1]) );
  INV_X1 U31 ( .A(n65), .ZN(Y[10]) );
  INV_X1 U32 ( .A(n37), .ZN(Y[7]) );
  INV_X1 U33 ( .A(n34), .ZN(Y[9]) );
  INV_X1 U34 ( .A(n43), .ZN(Y[30]) );
  AOI22_X1 U35 ( .A1(A[30]), .A2(SEL), .B1(B[30]), .B2(n69), .ZN(n43) );
  INV_X1 U36 ( .A(n49), .ZN(Y[25]) );
  AOI22_X1 U37 ( .A1(A[25]), .A2(SEL), .B1(B[25]), .B2(n70), .ZN(n49) );
  INV_X1 U38 ( .A(n46), .ZN(Y[28]) );
  AOI22_X1 U39 ( .A1(A[28]), .A2(SEL), .B1(B[28]), .B2(n69), .ZN(n46) );
  INV_X1 U40 ( .A(n53), .ZN(Y[21]) );
  AOI22_X1 U41 ( .A1(A[21]), .A2(SEL), .B1(B[21]), .B2(n71), .ZN(n53) );
  INV_X1 U42 ( .A(n50), .ZN(Y[24]) );
  AOI22_X1 U43 ( .A1(A[24]), .A2(SEL), .B1(B[24]), .B2(n70), .ZN(n50) );
  INV_X1 U44 ( .A(n47), .ZN(Y[27]) );
  AOI22_X1 U45 ( .A1(A[27]), .A2(SEL), .B1(B[27]), .B2(n70), .ZN(n47) );
  INV_X1 U46 ( .A(n62), .ZN(Y[13]) );
  INV_X1 U47 ( .A(n51), .ZN(Y[23]) );
  AOI22_X1 U48 ( .A1(A[23]), .A2(SEL), .B1(B[23]), .B2(n71), .ZN(n51) );
  INV_X1 U49 ( .A(n39), .ZN(Y[5]) );
  INV_X1 U50 ( .A(n45), .ZN(Y[29]) );
  AOI22_X1 U51 ( .A1(A[29]), .A2(SEL), .B1(B[29]), .B2(n69), .ZN(n45) );
  INV_X1 U52 ( .A(n54), .ZN(Y[20]) );
  AOI22_X1 U53 ( .A1(A[20]), .A2(SEL), .B1(B[20]), .B2(n71), .ZN(n54) );
  INV_X1 U54 ( .A(n56), .ZN(Y[19]) );
  AOI22_X1 U55 ( .A1(A[19]), .A2(SEL), .B1(B[19]), .B2(n72), .ZN(n56) );
  INV_X1 U56 ( .A(n60), .ZN(Y[15]) );
  AOI22_X1 U57 ( .A1(A[15]), .A2(SEL), .B1(B[15]), .B2(n73), .ZN(n60) );
  INV_X1 U58 ( .A(n66), .ZN(Y[0]) );
  AOI22_X1 U59 ( .A1(A[4]), .A2(SEL), .B1(B[4]), .B2(n68), .ZN(n40) );
  AOI22_X1 U60 ( .A1(A[3]), .A2(SEL), .B1(B[3]), .B2(n68), .ZN(n41) );
  AOI22_X1 U61 ( .A1(A[5]), .A2(SEL), .B1(B[5]), .B2(n68), .ZN(n39) );
  AOI22_X1 U62 ( .A1(A[6]), .A2(SEL), .B1(B[6]), .B2(n67), .ZN(n38) );
  AOI22_X1 U63 ( .A1(A[7]), .A2(SEL), .B1(B[7]), .B2(n67), .ZN(n37) );
  AOI22_X1 U64 ( .A1(A[8]), .A2(SEL), .B1(B[8]), .B2(n67), .ZN(n36) );
  AOI22_X1 U65 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n69), .ZN(n44) );
  AOI22_X1 U66 ( .A1(A[12]), .A2(SEL), .B1(B[12]), .B2(n74), .ZN(n63) );
  AOI22_X1 U67 ( .A1(A[13]), .A2(SEL), .B1(B[13]), .B2(n73), .ZN(n62) );
  AOI22_X1 U68 ( .A1(A[10]), .A2(SEL), .B1(B[10]), .B2(n74), .ZN(n65) );
  AOI22_X1 U69 ( .A1(A[11]), .A2(SEL), .B1(B[11]), .B2(n74), .ZN(n64) );
  AOI22_X1 U70 ( .A1(A[14]), .A2(SEL), .B1(B[14]), .B2(n73), .ZN(n61) );
  AOI22_X1 U71 ( .A1(SEL), .A2(A[9]), .B1(B[9]), .B2(n67), .ZN(n34) );
  AOI22_X1 U72 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n72), .ZN(n55) );
  AOI22_X1 U73 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n74), .ZN(n66) );
endmodule


module FD_INJ_NB5_1 ( CK, RESET, INJ_ZERO, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, INJ_ZERO;

  wire   [4:0] TMP_D;

  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U4 ( .A1(D[3]), .A2(INJ_ZERO), .ZN(TMP_D[3]) );
  AND2_X1 U5 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U6 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
  AND2_X1 U7 ( .A1(INJ_ZERO), .A2(D[4]), .ZN(TMP_D[4]) );
endmodule


module FD_INJ_NB5_2 ( CK, RESET, INJ_ZERO, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, INJ_ZERO;

  wire   [4:0] TMP_D;

  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U4 ( .A1(D[3]), .A2(INJ_ZERO), .ZN(TMP_D[3]) );
  AND2_X1 U5 ( .A1(INJ_ZERO), .A2(D[4]), .ZN(TMP_D[4]) );
  AND2_X1 U6 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U7 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
endmodule


module FD_INJ_NB5_0 ( CK, RESET, INJ_ZERO, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, INJ_ZERO;

  wire   [4:0] TMP_D;

  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[4]), .ZN(TMP_D[4]) );
  AND2_X1 U4 ( .A1(D[0]), .A2(INJ_ZERO), .ZN(TMP_D[0]) );
  AND2_X1 U5 ( .A1(D[1]), .A2(INJ_ZERO), .ZN(TMP_D[1]) );
  AND2_X1 U6 ( .A1(D[2]), .A2(INJ_ZERO), .ZN(TMP_D[2]) );
  AND2_X1 U7 ( .A1(D[3]), .A2(INJ_ZERO), .ZN(TMP_D[3]) );
endmodule


module MUX21_generic_NB5 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;
  wire   n7, n8, n9, n10, n11, n12;

  INV_X1 U1 ( .A(n7), .ZN(Y[4]) );
  AOI22_X1 U2 ( .A1(SEL), .A2(A[4]), .B1(B[4]), .B2(n8), .ZN(n7) );
  INV_X1 U3 ( .A(n12), .ZN(Y[0]) );
  AOI22_X1 U4 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n8), .ZN(n12) );
  INV_X1 U5 ( .A(n11), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n8), .ZN(n11) );
  INV_X1 U7 ( .A(n10), .ZN(Y[2]) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n8), .ZN(n10) );
  INV_X1 U9 ( .A(n9), .ZN(Y[3]) );
  AOI22_X1 U10 ( .A1(A[3]), .A2(SEL), .B1(B[3]), .B2(n8), .ZN(n9) );
  INV_X1 U11 ( .A(SEL), .ZN(n8) );
endmodule


module FD_INJ_NB32_2 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n38, n71, n72, n73, n74, n75, n76;
  wire   [31:0] TMP_D;
  assign n38 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n76), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n76), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n76), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n76), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n76), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n76), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n76), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n76), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n74), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n74), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n74), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n74), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n74), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n74), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n74), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n74), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n74), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n74), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n74), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n74), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n75), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n75), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n75), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n75), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n75), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n75), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n75), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n75), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n75), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n75), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n75), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n75), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n38), .Z(n75) );
  BUF_X1 U4 ( .A(n38), .Z(n74) );
  BUF_X1 U5 ( .A(n38), .Z(n76) );
  BUF_X1 U6 ( .A(INJ_ZERO), .Z(n71) );
  BUF_X1 U7 ( .A(INJ_ZERO), .Z(n72) );
  BUF_X1 U8 ( .A(INJ_ZERO), .Z(n73) );
  AND2_X1 U9 ( .A1(D[25]), .A2(n72), .ZN(TMP_D[25]) );
  AND2_X1 U10 ( .A1(D[26]), .A2(n72), .ZN(TMP_D[26]) );
  AND2_X1 U11 ( .A1(D[27]), .A2(n72), .ZN(TMP_D[27]) );
  AND2_X1 U12 ( .A1(D[28]), .A2(n72), .ZN(TMP_D[28]) );
  AND2_X1 U13 ( .A1(D[29]), .A2(n72), .ZN(TMP_D[29]) );
  AND2_X1 U14 ( .A1(D[30]), .A2(n72), .ZN(TMP_D[30]) );
  AND2_X1 U15 ( .A1(D[31]), .A2(n73), .ZN(TMP_D[31]) );
  AND2_X1 U16 ( .A1(D[0]), .A2(n71), .ZN(TMP_D[0]) );
  AND2_X1 U17 ( .A1(D[1]), .A2(n71), .ZN(TMP_D[1]) );
  AND2_X1 U18 ( .A1(D[2]), .A2(n72), .ZN(TMP_D[2]) );
  AND2_X1 U19 ( .A1(D[10]), .A2(n71), .ZN(TMP_D[10]) );
  AND2_X1 U20 ( .A1(D[11]), .A2(n71), .ZN(TMP_D[11]) );
  AND2_X1 U21 ( .A1(D[12]), .A2(n71), .ZN(TMP_D[12]) );
  AND2_X1 U22 ( .A1(D[13]), .A2(n71), .ZN(TMP_D[13]) );
  AND2_X1 U23 ( .A1(D[14]), .A2(n71), .ZN(TMP_D[14]) );
  AND2_X1 U24 ( .A1(D[15]), .A2(n71), .ZN(TMP_D[15]) );
  AND2_X1 U25 ( .A1(D[16]), .A2(n71), .ZN(TMP_D[16]) );
  AND2_X1 U26 ( .A1(D[17]), .A2(n71), .ZN(TMP_D[17]) );
  AND2_X1 U27 ( .A1(D[18]), .A2(n71), .ZN(TMP_D[18]) );
  AND2_X1 U28 ( .A1(D[19]), .A2(n71), .ZN(TMP_D[19]) );
  AND2_X1 U29 ( .A1(D[20]), .A2(n72), .ZN(TMP_D[20]) );
  AND2_X1 U30 ( .A1(D[21]), .A2(n72), .ZN(TMP_D[21]) );
  AND2_X1 U31 ( .A1(D[22]), .A2(n72), .ZN(TMP_D[22]) );
  AND2_X1 U32 ( .A1(D[23]), .A2(n72), .ZN(TMP_D[23]) );
  AND2_X1 U33 ( .A1(D[24]), .A2(n72), .ZN(TMP_D[24]) );
  AND2_X1 U34 ( .A1(n73), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U35 ( .A1(D[3]), .A2(n73), .ZN(TMP_D[3]) );
  AND2_X1 U36 ( .A1(D[4]), .A2(n73), .ZN(TMP_D[4]) );
  AND2_X1 U37 ( .A1(D[5]), .A2(n73), .ZN(TMP_D[5]) );
  AND2_X1 U38 ( .A1(D[6]), .A2(n73), .ZN(TMP_D[6]) );
  AND2_X1 U39 ( .A1(D[7]), .A2(n73), .ZN(TMP_D[7]) );
  AND2_X1 U40 ( .A1(D[8]), .A2(n73), .ZN(TMP_D[8]) );
endmodule


module SIGN_EXT_NB32 ( A, US, JMP, Y );
  input [25:0] A;
  output [31:0] Y;
  input US, JMP;
  wire   \Y[25] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  assign Y[31] = \Y[25] ;
  assign Y[30] = \Y[25] ;
  assign Y[29] = \Y[25] ;
  assign Y[28] = \Y[25] ;
  assign Y[27] = \Y[25] ;
  assign Y[26] = \Y[25] ;
  assign Y[25] = \Y[25] ;
  assign Y[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND2_X1 U2 ( .A1(n1), .A2(n11), .ZN(Y[16]) );
  NAND2_X1 U3 ( .A1(A[16]), .A2(JMP), .ZN(n11) );
  NAND2_X1 U4 ( .A1(n1), .A2(n10), .ZN(Y[17]) );
  NAND2_X1 U5 ( .A1(A[17]), .A2(JMP), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n1), .A2(n9), .ZN(Y[18]) );
  NAND2_X1 U7 ( .A1(A[18]), .A2(JMP), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n1), .A2(n8), .ZN(Y[19]) );
  NAND2_X1 U9 ( .A1(A[19]), .A2(JMP), .ZN(n8) );
  NAND2_X1 U10 ( .A1(n1), .A2(n7), .ZN(Y[20]) );
  NAND2_X1 U11 ( .A1(A[20]), .A2(JMP), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n1), .A2(n6), .ZN(Y[21]) );
  NAND2_X1 U13 ( .A1(A[21]), .A2(JMP), .ZN(n6) );
  NAND2_X1 U14 ( .A1(n1), .A2(n5), .ZN(Y[22]) );
  NAND2_X1 U15 ( .A1(A[22]), .A2(JMP), .ZN(n5) );
  NAND2_X1 U16 ( .A1(n1), .A2(n4), .ZN(Y[23]) );
  NAND2_X1 U17 ( .A1(A[23]), .A2(JMP), .ZN(n4) );
  NAND2_X1 U18 ( .A1(n1), .A2(n3), .ZN(Y[24]) );
  NAND2_X1 U19 ( .A1(A[24]), .A2(JMP), .ZN(n3) );
  NAND2_X1 U20 ( .A1(n12), .A2(\A[15] ), .ZN(n1) );
  NOR2_X1 U21 ( .A1(US), .A2(JMP), .ZN(n12) );
  NAND2_X1 U22 ( .A1(n1), .A2(n2), .ZN(\Y[25] ) );
  NAND2_X1 U23 ( .A1(JMP), .A2(A[25]), .ZN(n2) );
endmodule


module FD_INJ_NB32_3 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n38, n71, n72, n73, n74, n75, n76;
  wire   [31:0] TMP_D;
  assign n38 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n76), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n76), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n76), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n76), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n76), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n76), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n76), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n76), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n74), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n74), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n74), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n74), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n74), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n74), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n74), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n74), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n74), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n74), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n74), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n74), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n75), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n75), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n75), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n75), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n75), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n75), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n75), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n75), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n75), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n75), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n75), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n75), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n38), .Z(n75) );
  BUF_X1 U4 ( .A(n38), .Z(n74) );
  BUF_X1 U5 ( .A(n38), .Z(n76) );
  BUF_X1 U6 ( .A(INJ_ZERO), .Z(n71) );
  BUF_X1 U7 ( .A(INJ_ZERO), .Z(n72) );
  BUF_X1 U8 ( .A(INJ_ZERO), .Z(n73) );
  AND2_X1 U9 ( .A1(D[0]), .A2(n71), .ZN(TMP_D[0]) );
  AND2_X1 U10 ( .A1(D[1]), .A2(n71), .ZN(TMP_D[1]) );
  AND2_X1 U11 ( .A1(D[2]), .A2(n72), .ZN(TMP_D[2]) );
  AND2_X1 U12 ( .A1(D[10]), .A2(n71), .ZN(TMP_D[10]) );
  AND2_X1 U13 ( .A1(D[11]), .A2(n71), .ZN(TMP_D[11]) );
  AND2_X1 U14 ( .A1(D[12]), .A2(n71), .ZN(TMP_D[12]) );
  AND2_X1 U15 ( .A1(D[13]), .A2(n71), .ZN(TMP_D[13]) );
  AND2_X1 U16 ( .A1(D[14]), .A2(n71), .ZN(TMP_D[14]) );
  AND2_X1 U17 ( .A1(D[15]), .A2(n71), .ZN(TMP_D[15]) );
  AND2_X1 U18 ( .A1(D[16]), .A2(n71), .ZN(TMP_D[16]) );
  AND2_X1 U19 ( .A1(D[17]), .A2(n71), .ZN(TMP_D[17]) );
  AND2_X1 U20 ( .A1(D[18]), .A2(n71), .ZN(TMP_D[18]) );
  AND2_X1 U21 ( .A1(D[19]), .A2(n71), .ZN(TMP_D[19]) );
  AND2_X1 U22 ( .A1(D[20]), .A2(n72), .ZN(TMP_D[20]) );
  AND2_X1 U23 ( .A1(D[21]), .A2(n72), .ZN(TMP_D[21]) );
  AND2_X1 U24 ( .A1(D[22]), .A2(n72), .ZN(TMP_D[22]) );
  AND2_X1 U25 ( .A1(D[23]), .A2(n72), .ZN(TMP_D[23]) );
  AND2_X1 U26 ( .A1(D[24]), .A2(n72), .ZN(TMP_D[24]) );
  AND2_X1 U27 ( .A1(D[25]), .A2(n72), .ZN(TMP_D[25]) );
  AND2_X1 U28 ( .A1(D[26]), .A2(n72), .ZN(TMP_D[26]) );
  AND2_X1 U29 ( .A1(D[27]), .A2(n72), .ZN(TMP_D[27]) );
  AND2_X1 U30 ( .A1(D[28]), .A2(n72), .ZN(TMP_D[28]) );
  AND2_X1 U31 ( .A1(D[29]), .A2(n72), .ZN(TMP_D[29]) );
  AND2_X1 U32 ( .A1(D[30]), .A2(n72), .ZN(TMP_D[30]) );
  AND2_X1 U33 ( .A1(n73), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U34 ( .A1(D[3]), .A2(n73), .ZN(TMP_D[3]) );
  AND2_X1 U35 ( .A1(D[4]), .A2(n73), .ZN(TMP_D[4]) );
  AND2_X1 U36 ( .A1(D[5]), .A2(n73), .ZN(TMP_D[5]) );
  AND2_X1 U37 ( .A1(D[6]), .A2(n73), .ZN(TMP_D[6]) );
  AND2_X1 U38 ( .A1(D[7]), .A2(n73), .ZN(TMP_D[7]) );
  AND2_X1 U39 ( .A1(D[8]), .A2(n73), .ZN(TMP_D[8]) );
  AND2_X1 U40 ( .A1(D[31]), .A2(n73), .ZN(TMP_D[31]) );
endmodule


module FD_INJ_NB32_4 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n38, n71, n72, n73, n74, n75, n76;
  wire   [31:0] TMP_D;
  assign n38 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n76), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n76), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n76), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n76), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n76), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n76), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n76), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n76), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n74), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n74), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n74), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n74), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n74), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n74), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n74), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n74), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n74), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n74), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n74), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n74), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n75), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n75), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n75), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n75), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n75), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n75), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n75), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n75), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n75), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n75), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n75), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n75), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n38), .Z(n75) );
  BUF_X1 U4 ( .A(n38), .Z(n74) );
  BUF_X1 U5 ( .A(n38), .Z(n76) );
  AND2_X1 U6 ( .A1(D[1]), .A2(n71), .ZN(TMP_D[1]) );
  AND2_X1 U7 ( .A1(D[12]), .A2(n71), .ZN(TMP_D[12]) );
  AND2_X1 U8 ( .A1(D[13]), .A2(n71), .ZN(TMP_D[13]) );
  AND2_X1 U9 ( .A1(D[14]), .A2(n71), .ZN(TMP_D[14]) );
  AND2_X1 U10 ( .A1(D[15]), .A2(n71), .ZN(TMP_D[15]) );
  AND2_X1 U11 ( .A1(D[16]), .A2(n71), .ZN(TMP_D[16]) );
  AND2_X1 U12 ( .A1(D[17]), .A2(n71), .ZN(TMP_D[17]) );
  AND2_X1 U13 ( .A1(D[18]), .A2(n71), .ZN(TMP_D[18]) );
  AND2_X1 U14 ( .A1(D[19]), .A2(n71), .ZN(TMP_D[19]) );
  AND2_X1 U15 ( .A1(D[20]), .A2(n72), .ZN(TMP_D[20]) );
  AND2_X1 U16 ( .A1(D[21]), .A2(n72), .ZN(TMP_D[21]) );
  AND2_X1 U17 ( .A1(D[22]), .A2(n72), .ZN(TMP_D[22]) );
  AND2_X1 U18 ( .A1(D[23]), .A2(n72), .ZN(TMP_D[23]) );
  AND2_X1 U19 ( .A1(D[24]), .A2(n72), .ZN(TMP_D[24]) );
  AND2_X1 U20 ( .A1(D[25]), .A2(n72), .ZN(TMP_D[25]) );
  AND2_X1 U21 ( .A1(n73), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U22 ( .A1(D[4]), .A2(n73), .ZN(TMP_D[4]) );
  AND2_X1 U23 ( .A1(D[5]), .A2(n73), .ZN(TMP_D[5]) );
  AND2_X1 U24 ( .A1(D[6]), .A2(n73), .ZN(TMP_D[6]) );
  AND2_X1 U25 ( .A1(D[7]), .A2(n73), .ZN(TMP_D[7]) );
  AND2_X1 U26 ( .A1(D[8]), .A2(n73), .ZN(TMP_D[8]) );
  BUF_X1 U27 ( .A(INJ_ZERO), .Z(n71) );
  BUF_X1 U28 ( .A(INJ_ZERO), .Z(n72) );
  BUF_X1 U29 ( .A(INJ_ZERO), .Z(n73) );
  AND2_X1 U30 ( .A1(D[0]), .A2(n71), .ZN(TMP_D[0]) );
  AND2_X1 U31 ( .A1(D[2]), .A2(n72), .ZN(TMP_D[2]) );
  AND2_X1 U32 ( .A1(D[10]), .A2(n71), .ZN(TMP_D[10]) );
  AND2_X1 U33 ( .A1(D[11]), .A2(n71), .ZN(TMP_D[11]) );
  AND2_X1 U34 ( .A1(D[26]), .A2(n72), .ZN(TMP_D[26]) );
  AND2_X1 U35 ( .A1(D[27]), .A2(n72), .ZN(TMP_D[27]) );
  AND2_X1 U36 ( .A1(D[28]), .A2(n72), .ZN(TMP_D[28]) );
  AND2_X1 U37 ( .A1(D[29]), .A2(n72), .ZN(TMP_D[29]) );
  AND2_X1 U38 ( .A1(D[30]), .A2(n72), .ZN(TMP_D[30]) );
  AND2_X1 U39 ( .A1(D[3]), .A2(n73), .ZN(TMP_D[3]) );
  AND2_X1 U40 ( .A1(D[31]), .A2(n73), .ZN(TMP_D[31]) );
endmodule


module register_file_NB32_RS32 ( CLK, RESET, RD1, RD2, WR, ADD_WR, ADD_RD1, 
        ADD_RD2, DATAIN, HAZARD, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, RD1, RD2, WR;
  output HAZARD;
  wire   N4192, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n4, n5, n6, n7, n8, n9, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n3736, n3737, n3754, n3755, n3772,
         n3773, n3790, n3791, n3808, n3809, n3826, n3827, n3844, n3845, n3862,
         n3863, n3880, n3881, n3898, n3899, n3916, n3917, n3934, n3935, n3952,
         n3953, n3970, n3971, n3988, n3989, n4006, n4007, n4024, n4025, n4042,
         n4043, n4060, n4061, n4078, n4079, n4096, n4097, n4114, n4115, n4132,
         n4133, n4150, n4151, n4168, n4169, n4186, n4187, n4204, n4205, n4222,
         n4223, n4240, n4241, n4258, n4259, n4276, n4277, n4294, n4295,
         net86667, net86668, net86669, net86670, net86671, net86672, net86673,
         net86674, net86675, net86676, net86677, net86678, net86679, net86680,
         net86681, net86682, net86683, net86684, net86685, net86686, net86687,
         net86688, net86689, net86690, net86691, net86692, net86693, net86694,
         net86695, net86696, net86697, net86698, net86699, net86700, net86701,
         net86702, net86703, net86704, net86705, net86706, net86707, net86708,
         net86709, net86710, net86711, net86712, net86713, net86714, net86715,
         net86716, net86717, net86718, net86719, net86720, net86721, net86722,
         net86723, net86724, net86725, net86726, net86727, net86728, net86729,
         net86730, net86731, net86732, net86733, net86734, net86735, net86736,
         net86737, net86738, net86739, net86740, net86741, net86742, net86743,
         net86744, net86745, net86746, net86747, net86748, net86749, net86750,
         net86751, net86752, net86753, net86754, net86755, net86756, net86757,
         net86758, net86759, net86760, net86761, net86762, net86763, net86764,
         net86765, net86766, net86767, net86768, net86769, net86770, net86771,
         net86772, net86773, net86774, net86775, net86776, net86777, net86778,
         net86779, net86780, net86781, net86782, net86783, net86784, net86785,
         net86786, net86787, net86788, net86789, net86790, net86791, net86792,
         net86793, net86794, net86795, net86796, net86797, net86798, net86799,
         net86800, net86801, net86802, net86803, net86804, net86805, net86806,
         net86807, net86808, net86809, net86810, net86811, net86812, net86813,
         net86814, net86815, net86816, net86817, net86818, net86819, net86820,
         net86821, net86822, net86823, net86824, net86825, net86826, net86827,
         net86828, net86829, net86830, net86831, net86832, net86833, net86834,
         net86835, net86836, net86837, net86838, net86839, net86840, net86841,
         net86842, net86843, net86844, net86845, net86846, net86847, net86848,
         net86849, net86850, net86851, net86852, net86853, net86854, net86855,
         net86856, net86857, net86858, net86859, net86860, net86861, net86862,
         net86863, net86864, net86865, net86866, net86867, net86868, net86869,
         net86870, net86871, net86872, net86873, net86874, net86875, net86876,
         net86877, net86878, net86879, net86880, net86881, net86882, net86883,
         net86884, net86885, net86886, net86887, net86888, net86889, net86890,
         net86891, net86892, net86893, net86894, net86895, net86896, net86897,
         net86898, net86899, net86900, net86901, net86902, net86903, net86904,
         net86905, net86906, net86907, net86908, net86909, net86910, net86911,
         net86912, net86913, net86914, net86915, net86916, net86917, net86918,
         net86919, net86920, net86921, net86922, net86923, net86924, net86925,
         net86926, net86927, net86928, net86929, net86930, net86931, net86932,
         net86933, net86934, net86935, net86936, net86937, net86938, net86939,
         net86940, net86941, net86942, net86943, net86944, net86945, net86946,
         net86947, net86948, net86949, net86950, net86951, net86952, net86953,
         net86954, net86955, net86956, net86957, net86958, net86959, net86960,
         net86961, net86962, net86963, net86964, net86965, net86966, net86967,
         net86968, net86969, net86970, net86971, net86972, net86973, net86974,
         net86975, net86976, net86977, net86978, net86979, net86980, net86981,
         net86982, net86983, net86984, net86985, net86986, net86987, net86988,
         net86989, net86990, net86991, net86992, net86993, net86994, net86995,
         net86996, net86997, net86998, net86999, net87000, net87001, net87002,
         net87003, net87004, net87005, net87006, net87007, net87008, net87009,
         net87010, net87011, net87012, net87013, net87014, net87015, net87016,
         net87017, net87018, net87019, net87020, net87021, net87022, net87023,
         net87024, net87025, net87026, net87027, net87028, net87029, net87030,
         net87031, net87032, net87033, net87034, net87035, net87036, net87037,
         net87038, net87039, net87040, net87041, net87042, net87043, net87044,
         net87045, net87046, net87047, net87048, net87049, net87050, net87051,
         net87052, net87053, net87054, net87055, net87056, net87057, net87058,
         net87059, net87060, net87061, net87062, net87063, net87064, net87065,
         net87066, net87067, net87068, net87069, net87070, net87071, net87072,
         net87073, net87074, net87075, net87076, net87077, net87078, net87079,
         net87080, net87081, net87082, net87083, net87084, net87085, net87086,
         net87087, net87088, net87089, net87090, net87091, net87092, net87093,
         net87094, net87095, net87096, net87097, net87098, net87099, net87100,
         net87101, net87102, net87103, net87104, net87105, net87106, net87107,
         net87108, net87109, net87110, net87111, net87112, net87113, net87114,
         net87115, net87116, net87117, net87118, net87119, net87120, net87121,
         net87122, net87123, net87124, net87125, net87126, net87127, net87128,
         net87129, net87130, net87131, net87132, net87133, net87134, net87135,
         net87136, net87137, net87138, net87139, net87140, net87141, net87142,
         net87143, net87144, net87145, net87146, net87147, net87148, net87149,
         net87150, net87151, net87152, net87153, net87154, net87155, net87156,
         net87157, net87158, net87159, net87160, net87161, net87162, net87163,
         net87164, net87165, net87166, net87167, net87168, net87169, net87170,
         net87171, net87172, net87173, net87174, net87175, net87176, net87177,
         net87178, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1969, n1970, n1972, n1973, n1974, n1975, n1976, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2035, n2037, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2096,
         n2098, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2155, n2157, n2158, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2215, n2217, n2218, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2275, n2277, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2334, n2336, n2338, n2339, n2340, n2341, n2343, n2345, n2346,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736;

  DFF_X1 HAZARD_reg ( .D(N4192), .CK(CLK), .Q(HAZARD) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n3680), .CK(CLK), .QN(n1881) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n3679), .CK(CLK), .QN(n1883) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n3678), .CK(CLK), .QN(n1885) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n3677), .CK(CLK), .QN(n1887) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n3676), .CK(CLK), .QN(n1889) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n3675), .CK(CLK), .QN(n1891) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n3674), .CK(CLK), .QN(n1893) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n3673), .CK(CLK), .QN(n1895) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n3672), .CK(CLK), .QN(n1897) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n3671), .CK(CLK), .QN(n1899) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n3670), .CK(CLK), .QN(n1901) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n3669), .CK(CLK), .QN(n1903) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n3668), .CK(CLK), .QN(n1905) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n3667), .CK(CLK), .QN(n1907) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n3666), .CK(CLK), .QN(n1909) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n3665), .CK(CLK), .QN(n1911) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n3664), .CK(CLK), .QN(n1913) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n3663), .CK(CLK), .QN(n1915) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n3662), .CK(CLK), .QN(n1917) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n3661), .CK(CLK), .QN(n1919) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n3658), .CK(CLK), .QN(n1923) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n3657), .CK(CLK), .QN(n1925) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n3656), .CK(CLK), .QN(n1927) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n3655), .CK(CLK), .QN(n1929) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n3654), .CK(CLK), .QN(n1931) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n3653), .CK(CLK), .QN(n1933) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n3652), .CK(CLK), .QN(n1935) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n3651), .CK(CLK), .QN(n1937) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n3650), .CK(CLK), .QN(n1939) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n3641), .CK(CLK), .QN(n1945) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n3640), .CK(CLK), .QN(n1946) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n3639), .CK(CLK), .QN(n1947) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n3638), .CK(CLK), .QN(n1948) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n3637), .CK(CLK), .QN(n1949) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n3636), .CK(CLK), .QN(n1950) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n3635), .CK(CLK), .QN(n1951) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n3634), .CK(CLK), .QN(n1952) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n3633), .CK(CLK), .QN(n1953) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n3632), .CK(CLK), .QN(n1954) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n3631), .CK(CLK), .QN(n1955) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n3630), .CK(CLK), .QN(n1956) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n3629), .CK(CLK), .QN(n1957) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n3628), .CK(CLK), .QN(n1958) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n3627), .CK(CLK), .QN(n1959) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n3626), .CK(CLK), .QN(n1960) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n3624), .CK(CLK), .QN(n1961) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n3623), .CK(CLK), .QN(n1962) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n3622), .CK(CLK), .QN(n1963) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n3621), .CK(CLK), .QN(n1964) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n3618), .CK(CLK), .QN(n1965) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n3617), .CK(CLK), .QN(n1966) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n3552), .CK(CLK), .QN(n1979) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n3551), .CK(CLK), .QN(n1980) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n3550), .CK(CLK), .QN(n1981) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n3549), .CK(CLK), .QN(n1982) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n3548), .CK(CLK), .QN(n1983) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n3547), .CK(CLK), .QN(n1984) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n3546), .CK(CLK), .QN(n1985) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n3545), .CK(CLK), .QN(n1986) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n3544), .CK(CLK), .QN(n1987) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n3543), .CK(CLK), .QN(n1988) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n3542), .CK(CLK), .QN(n1989) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n3541), .CK(CLK), .QN(n1990) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n3540), .CK(CLK), .QN(n1991) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n3539), .CK(CLK), .QN(n1992) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n3538), .CK(CLK), .QN(n1993) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n3537), .CK(CLK), .QN(n1994) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n3536), .CK(CLK), .QN(n1995) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n3535), .CK(CLK), .QN(n1996) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n3534), .CK(CLK), .QN(n1997) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n3533), .CK(CLK), .QN(n1998) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n3530), .CK(CLK), .QN(n1999) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n3529), .CK(CLK), .QN(n2000) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n3528), .CK(CLK), .QN(n2001) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n3527), .CK(CLK), .QN(n2002) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n3526), .CK(CLK), .QN(n2003) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n3525), .CK(CLK), .QN(n2004) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n3524), .CK(CLK), .QN(n2005) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n3523), .CK(CLK), .QN(n2006) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n3522), .CK(CLK), .QN(n2007) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n3514), .CK(CLK), .QN(n2011) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n3513), .CK(CLK), .QN(n2012) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n3512), .CK(CLK), .QN(n2013) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n3511), .CK(CLK), .QN(n2014) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n3510), .CK(CLK), .QN(n2015) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n3509), .CK(CLK), .QN(n2016) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n3508), .CK(CLK), .QN(n2017) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n3507), .CK(CLK), .QN(n2018) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n3506), .CK(CLK), .QN(n2019) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n3505), .CK(CLK), .QN(n2020) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n3504), .CK(CLK), .QN(n2021) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n3503), .CK(CLK), .QN(n2022) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n3502), .CK(CLK), .QN(n2023) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n3501), .CK(CLK), .QN(n2024) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n3500), .CK(CLK), .QN(n2025) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n3499), .CK(CLK), .QN(n2026) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n3498), .CK(CLK), .QN(n2027) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n3496), .CK(CLK), .QN(n2028) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n3495), .CK(CLK), .QN(n2029) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n3494), .CK(CLK), .QN(n2030) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n3493), .CK(CLK), .QN(n2031) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n3490), .CK(CLK), .QN(n2032) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n3489), .CK(CLK), .QN(n2033) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n3424), .CK(CLK), .QN(n2040) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n3423), .CK(CLK), .QN(n2041) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n3422), .CK(CLK), .QN(n2042) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n3421), .CK(CLK), .QN(n2043) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n3420), .CK(CLK), .QN(n2044) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n3419), .CK(CLK), .QN(n2045) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n3418), .CK(CLK), .QN(n2046) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n3417), .CK(CLK), .QN(n2047) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n3416), .CK(CLK), .QN(n2048) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n3415), .CK(CLK), .QN(n2049) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n3414), .CK(CLK), .QN(n2050) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n3413), .CK(CLK), .QN(n2051) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n3412), .CK(CLK), .QN(n2052) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n3411), .CK(CLK), .QN(n2053) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n3410), .CK(CLK), .QN(n2054) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n3409), .CK(CLK), .QN(n2055) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n3408), .CK(CLK), .QN(n2056) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n3407), .CK(CLK), .QN(n2057) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n3406), .CK(CLK), .QN(n2058) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n3402), .CK(CLK), .QN(n2059) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n3401), .CK(CLK), .QN(n2060) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n3400), .CK(CLK), .QN(n2061) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n3399), .CK(CLK), .QN(n2062) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n3398), .CK(CLK), .QN(n2063) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n3397), .CK(CLK), .QN(n2064) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n3396), .CK(CLK), .QN(n2065) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n3395), .CK(CLK), .QN(n2066) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n3394), .CK(CLK), .QN(n2067) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n3386), .CK(CLK), .QN(n2071) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n3385), .CK(CLK), .QN(n2072) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n3384), .CK(CLK), .QN(n2073) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n3383), .CK(CLK), .QN(n2074) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n3382), .CK(CLK), .QN(n2075) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n3381), .CK(CLK), .QN(n2076) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n3380), .CK(CLK), .QN(n2077) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n3379), .CK(CLK), .QN(n2078) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n3378), .CK(CLK), .QN(n2079) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n3377), .CK(CLK), .QN(n2080) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n3376), .CK(CLK), .QN(n2081) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n3375), .CK(CLK), .QN(n2082) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n3374), .CK(CLK), .QN(n2083) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n3373), .CK(CLK), .QN(n2084) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n3372), .CK(CLK), .QN(n2085) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n3371), .CK(CLK), .QN(n2086) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n3370), .CK(CLK), .QN(n2087) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n3369), .CK(CLK), .QN(n2088) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n3368), .CK(CLK), .QN(n2089) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n3367), .CK(CLK), .QN(n2090) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n3366), .CK(CLK), .QN(n2091) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n3365), .CK(CLK), .QN(n2092) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n3362), .CK(CLK), .QN(n2093) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n3361), .CK(CLK), .QN(n2094) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n3296), .CK(CLK), .QN(n2101) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n3295), .CK(CLK), .QN(n2102) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n3294), .CK(CLK), .QN(n2103) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n3293), .CK(CLK), .QN(n2104) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n3292), .CK(CLK), .QN(n2105) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n3291), .CK(CLK), .QN(n2106) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n3290), .CK(CLK), .QN(n2107) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n3289), .CK(CLK), .QN(n2108) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n3288), .CK(CLK), .QN(n2109) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n3287), .CK(CLK), .QN(n2110) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n3286), .CK(CLK), .QN(n2111) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n3285), .CK(CLK), .QN(n2112) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n3284), .CK(CLK), .QN(n2113) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n3283), .CK(CLK), .QN(n2114) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n3282), .CK(CLK), .QN(n2115) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n3281), .CK(CLK), .QN(n2116) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n3280), .CK(CLK), .QN(n2117) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n3279), .CK(CLK), .QN(n2118) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n3278), .CK(CLK), .QN(n2119) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n3274), .CK(CLK), .QN(n2120) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n3273), .CK(CLK), .QN(n2121) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n3272), .CK(CLK), .QN(n2122) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n3271), .CK(CLK), .QN(n2123) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n3270), .CK(CLK), .QN(n2124) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n3269), .CK(CLK), .QN(n2125) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n3268), .CK(CLK), .QN(n2126) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n3267), .CK(CLK), .QN(n2127) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n3266), .CK(CLK), .QN(n2128) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n3258), .CK(CLK), .QN(n2132) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n3257), .CK(CLK), .QN(n2133) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n3256), .CK(CLK), .QN(n2134) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n3255), .CK(CLK), .QN(n2135) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n3254), .CK(CLK), .QN(n2136) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n3253), .CK(CLK), .QN(n2137) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n3252), .CK(CLK), .QN(n2138) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n3251), .CK(CLK), .QN(n2139) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n3250), .CK(CLK), .QN(n2140) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n3249), .CK(CLK), .QN(n2141) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n3248), .CK(CLK), .QN(n2142) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n3247), .CK(CLK), .QN(n2143) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n3246), .CK(CLK), .QN(n2144) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n3245), .CK(CLK), .QN(n2145) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n3244), .CK(CLK), .QN(n2146) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n3243), .CK(CLK), .QN(n2147) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n3241), .CK(CLK), .QN(n2148) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n3240), .CK(CLK), .QN(n2149) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n3239), .CK(CLK), .QN(n2150) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n3238), .CK(CLK), .QN(n2151) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n3234), .CK(CLK), .QN(n2152) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n3233), .CK(CLK), .QN(n2153) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n3162), .CK(CLK), .QN(n2161) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n3161), .CK(CLK), .QN(n2162) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n3160), .CK(CLK), .QN(n2163) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n3159), .CK(CLK), .QN(n2164) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n3158), .CK(CLK), .QN(n2165) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n3157), .CK(CLK), .QN(n2166) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n3156), .CK(CLK), .QN(n2167) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n3155), .CK(CLK), .QN(n2168) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n3154), .CK(CLK), .QN(n2169) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n3153), .CK(CLK), .QN(n2170) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n3152), .CK(CLK), .QN(n2171) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n3151), .CK(CLK), .QN(n2172) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n3150), .CK(CLK), .QN(n2173) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n3149), .CK(CLK), .QN(n2174) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n3148), .CK(CLK), .QN(n2175) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n3147), .CK(CLK), .QN(n2176) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n3145), .CK(CLK), .QN(n2177) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n3144), .CK(CLK), .QN(n2178) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n3143), .CK(CLK), .QN(n2179) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n3142), .CK(CLK), .QN(n2180) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n3138), .CK(CLK), .QN(n2181) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n3137), .CK(CLK), .QN(n2182) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n3136), .CK(CLK), .QN(n2186) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n3135), .CK(CLK), .QN(n2187) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n3134), .CK(CLK), .QN(n2188) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n3133), .CK(CLK), .QN(n2189) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n3132), .CK(CLK), .QN(n2190) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n3131), .CK(CLK), .QN(n2191) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n3130), .CK(CLK), .QN(n2192) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n3129), .CK(CLK), .QN(n2193) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n3128), .CK(CLK), .QN(n2194) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n3127), .CK(CLK), .QN(n2195) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n3126), .CK(CLK), .QN(n2196) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n3125), .CK(CLK), .QN(n2197) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n3124), .CK(CLK), .QN(n2198) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n3123), .CK(CLK), .QN(n2199) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n3122), .CK(CLK), .QN(n2200) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n3121), .CK(CLK), .QN(n2201) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n3120), .CK(CLK), .QN(n2202) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n3119), .CK(CLK), .QN(n2203) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n3118), .CK(CLK), .QN(n2204) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n3114), .CK(CLK), .QN(n2205) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n3113), .CK(CLK), .QN(n2206) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n3112), .CK(CLK), .QN(n2207) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n3111), .CK(CLK), .QN(n2208) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n3110), .CK(CLK), .QN(n2209) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n3109), .CK(CLK), .QN(n2210) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n3108), .CK(CLK), .QN(n2211) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n3107), .CK(CLK), .QN(n2212) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n3106), .CK(CLK), .QN(n2213) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n3034), .CK(CLK), .QN(n2221) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n3033), .CK(CLK), .QN(n2222) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n3032), .CK(CLK), .QN(n2223) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n3031), .CK(CLK), .QN(n2224) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n3030), .CK(CLK), .QN(n2225) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n3029), .CK(CLK), .QN(n2226) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n3028), .CK(CLK), .QN(n2227) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n3027), .CK(CLK), .QN(n2228) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n3026), .CK(CLK), .QN(n2229) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n3025), .CK(CLK), .QN(n2230) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n3024), .CK(CLK), .QN(n2231) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n3023), .CK(CLK), .QN(n2232) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n3022), .CK(CLK), .QN(n2233) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n3021), .CK(CLK), .QN(n2234) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n3020), .CK(CLK), .QN(n2235) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n3019), .CK(CLK), .QN(n2236) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n3017), .CK(CLK), .QN(n2237) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n3016), .CK(CLK), .QN(n2238) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n3015), .CK(CLK), .QN(n2239) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n3014), .CK(CLK), .QN(n2240) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n3010), .CK(CLK), .QN(n2241) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n3009), .CK(CLK), .QN(n2242) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n3008), .CK(CLK), .QN(n2246) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n3007), .CK(CLK), .QN(n2247) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n3006), .CK(CLK), .QN(n2248) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n3005), .CK(CLK), .QN(n2249) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n3004), .CK(CLK), .QN(n2250) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n3003), .CK(CLK), .QN(n2251) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n3002), .CK(CLK), .QN(n2252) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n3001), .CK(CLK), .QN(n2253) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n3000), .CK(CLK), .QN(n2254) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n2999), .CK(CLK), .QN(n2255) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n2998), .CK(CLK), .QN(n2256) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n2997), .CK(CLK), .QN(n2257) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n2996), .CK(CLK), .QN(n2258) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n2995), .CK(CLK), .QN(n2259) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n2994), .CK(CLK), .QN(n2260) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n2993), .CK(CLK), .QN(n2261) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n2992), .CK(CLK), .QN(n2262) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n2991), .CK(CLK), .QN(n2263) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n2990), .CK(CLK), .QN(n2264) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n2986), .CK(CLK), .QN(n2265) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n2985), .CK(CLK), .QN(n2266) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n2984), .CK(CLK), .QN(n2267) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n2983), .CK(CLK), .QN(n2268) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n2982), .CK(CLK), .QN(n2269) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n2981), .CK(CLK), .QN(n2270) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n2980), .CK(CLK), .QN(n2271) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n2979), .CK(CLK), .QN(n2272) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n2978), .CK(CLK), .QN(n2273) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n2912), .CK(CLK), .QN(n2280) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n2911), .CK(CLK), .QN(n2281) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n2910), .CK(CLK), .QN(n2282) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n2909), .CK(CLK), .QN(n2283) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n2908), .CK(CLK), .QN(n2284) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n2907), .CK(CLK), .QN(n2285) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n2906), .CK(CLK), .QN(n2286) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n2905), .CK(CLK), .QN(n2287) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n2904), .CK(CLK), .QN(n2288) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n2903), .CK(CLK), .QN(n2289) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n2902), .CK(CLK), .QN(n2290) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n2901), .CK(CLK), .QN(n2291) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n2900), .CK(CLK), .QN(n2292) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n2899), .CK(CLK), .QN(n2293) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n2898), .CK(CLK), .QN(n2294) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n2897), .CK(CLK), .QN(n2295) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n2896), .CK(CLK), .QN(n2296) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n2895), .CK(CLK), .QN(n2297) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n2894), .CK(CLK), .QN(n2298) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n2890), .CK(CLK), .QN(n2299) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n2889), .CK(CLK), .QN(n2300) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n2888), .CK(CLK), .QN(n2301) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n2887), .CK(CLK), .QN(n2302) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n2886), .CK(CLK), .QN(n2303) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n2885), .CK(CLK), .QN(n2304) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n2884), .CK(CLK), .QN(n2305) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n2883), .CK(CLK), .QN(n2306) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n2882), .CK(CLK), .QN(n2307) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n2874), .CK(CLK), .QN(n2311) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n2873), .CK(CLK), .QN(n2312) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n2872), .CK(CLK), .QN(n2313) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n2871), .CK(CLK), .QN(n2314) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n2870), .CK(CLK), .QN(n2315) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n2869), .CK(CLK), .QN(n2316) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n2868), .CK(CLK), .QN(n2317) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n2867), .CK(CLK), .QN(n2318) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n2866), .CK(CLK), .QN(n2319) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n2865), .CK(CLK), .QN(n2320) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n2864), .CK(CLK), .QN(n2321) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n2863), .CK(CLK), .QN(n2322) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n2862), .CK(CLK), .QN(n2323) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n2861), .CK(CLK), .QN(n2324) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n2860), .CK(CLK), .QN(n2325) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n2859), .CK(CLK), .QN(n2326) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n2857), .CK(CLK), .QN(n2327) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n2856), .CK(CLK), .QN(n2328) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n2855), .CK(CLK), .QN(n2329) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n2854), .CK(CLK), .QN(n2330) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n2850), .CK(CLK), .QN(n2331) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n2849), .CK(CLK), .QN(n2332) );
  NOR3_X2 U1770 ( .A1(n5081), .A2(ADD_RD2[2]), .A3(n5082), .ZN(n5051) );
  NOR3_X2 U1773 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n5082), .ZN(n5052) );
  NOR3_X2 U1778 ( .A1(n5082), .A2(n5081), .A3(n5086), .ZN(n5045) );
  NOR3_X2 U1783 ( .A1(n5082), .A2(ADD_RD2[1]), .A3(n5086), .ZN(n5047) );
  NOR3_X2 U3290 ( .A1(n5709), .A2(ADD_RD1[2]), .A3(n5710), .ZN(n5689) );
  NOR3_X2 U3294 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n5710), .ZN(n5690) );
  NOR3_X2 U3301 ( .A1(n5710), .A2(n5709), .A3(n5712), .ZN(n5685) );
  NOR3_X2 U3306 ( .A1(n5710), .A2(ADD_RD1[1]), .A3(n5712), .ZN(n5687) );
  NAND3_X1 U3333 ( .A1(n1974), .A2(n1975), .A3(n1976), .ZN(n1941) );
  NAND3_X1 U3334 ( .A1(n1976), .A2(n1975), .A3(ADD_WR[2]), .ZN(n2008) );
  NAND3_X1 U3335 ( .A1(n1976), .A2(n1974), .A3(ADD_WR[3]), .ZN(n2068) );
  NAND3_X1 U3336 ( .A1(ADD_WR[2]), .A2(n1976), .A3(ADD_WR[3]), .ZN(n2129) );
  NAND3_X1 U3337 ( .A1(n1974), .A2(n1975), .A3(n2218), .ZN(n2183) );
  NAND3_X1 U3338 ( .A1(ADD_WR[2]), .A2(n1975), .A3(n2218), .ZN(n2243) );
  NAND3_X1 U3339 ( .A1(ADD_WR[3]), .A2(n1974), .A3(n2218), .ZN(n2308) );
  NAND3_X1 U3340 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .A3(n2218), .ZN(n2339) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n2664), .CK(CLK), .Q(n2481), .QN(net86674) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2663), .CK(CLK), .Q(n2515), .QN(net86673) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2662), .CK(CLK), .Q(n2549), .QN(net86672) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n2661), .CK(CLK), .Q(n2583), .QN(net86671) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2660), .CK(CLK), .Q(n2617), .QN(net86670) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n2659), .CK(CLK), .Q(n4320), .QN(net86669) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n2658), .CK(CLK), .Q(n4694), .QN(net86668) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n2657), .CK(CLK), .Q(n5085), .QN(net86667) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n2688), .CK(CLK), .Q(n2651), .QN(
        net86698) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n2687), .CK(CLK), .Q(n3710), .QN(
        net86697) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2686), .CK(CLK), .Q(n4354), .QN(
        net86696) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n2685), .CK(CLK), .Q(n4388), .QN(
        net86695) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n2684), .CK(CLK), .Q(n4422), .QN(
        net86694) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2683), .CK(CLK), .Q(n4456), .QN(
        net86693) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n2682), .CK(CLK), .Q(n4490), .QN(
        net86692) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2681), .CK(CLK), .Q(n4524), .QN(
        net86691) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n2680), .CK(CLK), .Q(n4558), .QN(
        net86690) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2679), .CK(CLK), .Q(n4592), .QN(
        net86689) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n2678), .CK(CLK), .Q(n4626), .QN(
        net86688) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2677), .CK(CLK), .Q(n4660), .QN(
        net86687) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n2676), .CK(CLK), .Q(n4728), .QN(
        net86686) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n2675), .CK(CLK), .Q(n4762), .QN(
        net86685) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n2674), .CK(CLK), .Q(n4796), .QN(
        net86684) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n2673), .CK(CLK), .Q(n4830), .QN(
        net86683) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n2672), .CK(CLK), .Q(n4864), .QN(
        net86682) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n2671), .CK(CLK), .Q(n4898), .QN(
        net86681) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n2670), .CK(CLK), .Q(n4932), .QN(
        net86680) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n2669), .CK(CLK), .Q(n4966), .QN(
        net86679) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n2668), .CK(CLK), .Q(n5000), .QN(
        net86678) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2667), .CK(CLK), .Q(n5034), .QN(
        net86677) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n2666), .CK(CLK), .Q(n2413), .QN(net86676) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n2665), .CK(CLK), .Q(n2447), .QN(net86675) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n3648), .CK(CLK), .QN(n50) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n3647), .CK(CLK), .QN(n57) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n3646), .CK(CLK), .QN(n71) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n3645), .CK(CLK), .QN(n78) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n3644), .CK(CLK), .QN(n85) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n3643), .CK(CLK), .QN(n92) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n3642), .CK(CLK), .QN(n99) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n3625), .CK(CLK), .QN(n8) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n3620), .CK(CLK), .QN(n43) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n3619), .CK(CLK), .QN(n64) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n2720), .CK(CLK), .Q(n2650), .QN(
        net86730) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n2719), .CK(CLK), .Q(n3709), .QN(
        net86729) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2718), .CK(CLK), .Q(n4353), .QN(
        net86728) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2717), .CK(CLK), .Q(n4387), .QN(
        net86727) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n2716), .CK(CLK), .Q(n4421), .QN(
        net86726) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2715), .CK(CLK), .Q(n4455), .QN(
        net86725) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n2714), .CK(CLK), .Q(n4489), .QN(
        net86724) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n2713), .CK(CLK), .Q(n4523), .QN(
        net86723) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n2784), .CK(CLK), .QN(n3862) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n2783), .CK(CLK), .QN(n3880) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n2782), .CK(CLK), .QN(n3916) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n2781), .CK(CLK), .QN(n3934) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n2780), .CK(CLK), .QN(n3952) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n2779), .CK(CLK), .QN(n3970) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n2778), .CK(CLK), .QN(n3988) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n2777), .CK(CLK), .QN(n4006) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n2752), .CK(CLK), .QN(n3863) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n2751), .CK(CLK), .QN(n3881) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n2750), .CK(CLK), .QN(n3917) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n2749), .CK(CLK), .QN(n3935) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n2748), .CK(CLK), .QN(n3953) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n2747), .CK(CLK), .QN(n3971) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n2746), .CK(CLK), .QN(n3989) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n2745), .CK(CLK), .QN(n4007) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n2816), .CK(CLK), .Q(n2647), .QN(
        net86762) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n2815), .CK(CLK), .Q(n3706), .QN(
        net86761) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2814), .CK(CLK), .Q(n4350), .QN(
        net86760) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2813), .CK(CLK), .Q(n4384), .QN(
        net86759) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n2812), .CK(CLK), .Q(n4418), .QN(
        net86758) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2811), .CK(CLK), .Q(n4452), .QN(
        net86757) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n2810), .CK(CLK), .Q(n4486), .QN(
        net86756) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2809), .CK(CLK), .Q(n4520), .QN(
        net86755) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n2848), .CK(CLK), .Q(n2648), .QN(
        net86794) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n2847), .CK(CLK), .Q(n3707), .QN(
        net86793) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n2846), .CK(CLK), .Q(n4351), .QN(
        net86792) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n2845), .CK(CLK), .Q(n4385), .QN(
        net86791) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n2844), .CK(CLK), .Q(n4419), .QN(
        net86790) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n2843), .CK(CLK), .Q(n4453), .QN(
        net86789) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n2842), .CK(CLK), .Q(n4487), .QN(
        net86788) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n2841), .CK(CLK), .Q(n4521), .QN(
        net86787) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n2944), .CK(CLK), .Q(n2641), .QN(
        net86826) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n2943), .CK(CLK), .Q(n3700), .QN(
        net86825) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n2942), .CK(CLK), .Q(n4344), .QN(
        net86824) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n2941), .CK(CLK), .Q(n4378), .QN(
        net86823) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n2940), .CK(CLK), .Q(n4412), .QN(
        net86822) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n2939), .CK(CLK), .Q(n4446), .QN(
        net86821) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n2938), .CK(CLK), .Q(n4480), .QN(
        net86820) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n2937), .CK(CLK), .Q(n4514), .QN(
        net86819) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n2976), .CK(CLK), .Q(n2642), .QN(
        net86858) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n2975), .CK(CLK), .Q(n3701), .QN(
        net86857) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n2974), .CK(CLK), .Q(n4345), .QN(
        net86856) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n2973), .CK(CLK), .Q(n4379), .QN(
        net86855) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n2972), .CK(CLK), .Q(n4413), .QN(
        net86854) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n2971), .CK(CLK), .Q(n4447), .QN(
        net86853) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n2970), .CK(CLK), .Q(n4481), .QN(
        net86852) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n2969), .CK(CLK), .Q(n4515), .QN(
        net86851) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n3072), .CK(CLK), .Q(n2644), .QN(
        net86890) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n3071), .CK(CLK), .Q(n3703), .QN(
        net86889) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n3070), .CK(CLK), .Q(n4347), .QN(
        net86888) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n3069), .CK(CLK), .Q(n4381), .QN(
        net86887) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n3068), .CK(CLK), .Q(n4415), .QN(
        net86886) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n3067), .CK(CLK), .Q(n4449), .QN(
        net86885) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n3066), .CK(CLK), .Q(n4483), .QN(
        net86884) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n3065), .CK(CLK), .Q(n4517), .QN(
        net86883) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n3104), .CK(CLK), .Q(n2645), .QN(
        net86922) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n3103), .CK(CLK), .Q(n3704), .QN(
        net86921) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n3102), .CK(CLK), .Q(n4348), .QN(
        net86920) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n3101), .CK(CLK), .Q(n4382), .QN(
        net86919) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n3100), .CK(CLK), .Q(n4416), .QN(
        net86918) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n3099), .CK(CLK), .Q(n4450), .QN(
        net86917) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n3098), .CK(CLK), .Q(n4484), .QN(
        net86916) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n3097), .CK(CLK), .Q(n4518), .QN(
        net86915) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n3200), .CK(CLK), .Q(n2626), .QN(
        net86954) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n3199), .CK(CLK), .Q(n3685), .QN(
        net86953) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n3198), .CK(CLK), .Q(n4329), .QN(
        net86952) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n3197), .CK(CLK), .Q(n4363), .QN(
        net86951) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n3196), .CK(CLK), .Q(n4397), .QN(
        net86950) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n3195), .CK(CLK), .Q(n4431), .QN(
        net86949) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n3194), .CK(CLK), .Q(n4465), .QN(
        net86948) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n3193), .CK(CLK), .Q(n4499), .QN(
        net86947) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n3232), .CK(CLK), .Q(n2625), .QN(
        net86986) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n3231), .CK(CLK), .Q(n3684), .QN(
        net86985) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n3230), .CK(CLK), .Q(n4328), .QN(
        net86984) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n3229), .CK(CLK), .Q(n4362), .QN(
        net86983) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n3228), .CK(CLK), .Q(n4396), .QN(
        net86982) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n3227), .CK(CLK), .Q(n4430), .QN(
        net86981) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n3226), .CK(CLK), .Q(n4464), .QN(
        net86980) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n3225), .CK(CLK), .Q(n4498), .QN(
        net86979) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n3328), .CK(CLK), .Q(n2629), .QN(
        net87018) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n3327), .CK(CLK), .Q(n3688), .QN(
        net87017) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n3326), .CK(CLK), .Q(n4332), .QN(
        net87016) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n3325), .CK(CLK), .Q(n4366), .QN(
        net87015) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n3324), .CK(CLK), .Q(n4400), .QN(
        net87014) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n3323), .CK(CLK), .Q(n4434), .QN(
        net87013) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n3322), .CK(CLK), .Q(n4468), .QN(
        net87012) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n3321), .CK(CLK), .Q(n4502), .QN(
        net87011) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n3360), .CK(CLK), .Q(n2628), .QN(
        net87050) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n3359), .CK(CLK), .Q(n3687), .QN(
        net87049) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n3358), .CK(CLK), .Q(n4331), .QN(
        net87048) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n3357), .CK(CLK), .Q(n4365), .QN(
        net87047) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n3356), .CK(CLK), .Q(n4399), .QN(
        net87046) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n3355), .CK(CLK), .Q(n4433), .QN(
        net87045) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n3354), .CK(CLK), .Q(n4467), .QN(
        net87044) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n3353), .CK(CLK), .Q(n4501), .QN(
        net87043) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n3456), .CK(CLK), .Q(n2632), .QN(net87082) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n3455), .CK(CLK), .Q(n3691), .QN(net87081) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n3454), .CK(CLK), .Q(n4335), .QN(net87080) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n3453), .CK(CLK), .Q(n4369), .QN(net87079) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n3452), .CK(CLK), .Q(n4403), .QN(net87078) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n3451), .CK(CLK), .Q(n4437), .QN(net87077) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n3450), .CK(CLK), .Q(n4471), .QN(net87076) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n3449), .CK(CLK), .Q(n4505), .QN(net87075) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n3488), .CK(CLK), .Q(n2631), .QN(net87114) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n3487), .CK(CLK), .Q(n3690), .QN(net87113) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n3486), .CK(CLK), .Q(n4334), .QN(net87112) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n3485), .CK(CLK), .Q(n4368), .QN(net87111) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n3484), .CK(CLK), .Q(n4402), .QN(net87110) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n3483), .CK(CLK), .Q(n4436), .QN(net87109) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n3482), .CK(CLK), .Q(n4470), .QN(net87108) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n3481), .CK(CLK), .Q(n4504), .QN(net87107) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n3616), .CK(CLK), .Q(n2634), .QN(net87178) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n3615), .CK(CLK), .Q(n3693), .QN(net87177) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n3614), .CK(CLK), .Q(n4337), .QN(net87176) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n3613), .CK(CLK), .Q(n4371), .QN(net87175) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n3612), .CK(CLK), .Q(n4405), .QN(net87174) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n3611), .CK(CLK), .Q(n4439), .QN(net87173) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n3610), .CK(CLK), .Q(n4473), .QN(net87172) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n3609), .CK(CLK), .Q(n4507), .QN(net87171) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n3584), .CK(CLK), .Q(n2635), .QN(net87146) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n3583), .CK(CLK), .Q(n3694), .QN(net87145) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n3582), .CK(CLK), .Q(n4338), .QN(net87144) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n3581), .CK(CLK), .Q(n4372), .QN(net87143) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n3580), .CK(CLK), .Q(n4406), .QN(net87142) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n3579), .CK(CLK), .Q(n4440), .QN(net87141) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n3578), .CK(CLK), .Q(n4474), .QN(net87140) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n3577), .CK(CLK), .Q(n4508), .QN(net87139) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n2712), .CK(CLK), .Q(n4557), .QN(
        net86722) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2711), .CK(CLK), .Q(n4591), .QN(
        net86721) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n2710), .CK(CLK), .Q(n4625), .QN(
        net86720) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2709), .CK(CLK), .Q(n4659), .QN(
        net86719) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n2708), .CK(CLK), .Q(n4727), .QN(
        net86718) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n2707), .CK(CLK), .Q(n4761), .QN(
        net86717) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n2706), .CK(CLK), .Q(n4795), .QN(
        net86716) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n2705), .CK(CLK), .Q(n4829), .QN(
        net86715) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n2704), .CK(CLK), .Q(n4863), .QN(
        net86714) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n2703), .CK(CLK), .Q(n4897), .QN(
        net86713) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n2702), .CK(CLK), .Q(n4931), .QN(
        net86712) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n2701), .CK(CLK), .Q(n4965), .QN(
        net86711) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n2700), .CK(CLK), .Q(n4999), .QN(
        net86710) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2699), .CK(CLK), .Q(n5033), .QN(
        net86709) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n2698), .CK(CLK), .Q(n2411), .QN(net86708) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n2697), .CK(CLK), .Q(n2446), .QN(net86707) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n2696), .CK(CLK), .Q(n2480), .QN(net86706) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2695), .CK(CLK), .Q(n2514), .QN(net86705) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2694), .CK(CLK), .Q(n2548), .QN(net86704) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n2693), .CK(CLK), .Q(n2582), .QN(net86703) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2692), .CK(CLK), .Q(n2616), .QN(net86702) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n2691), .CK(CLK), .Q(n4319), .QN(net86701) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n2690), .CK(CLK), .Q(n4693), .QN(net86700) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n2689), .CK(CLK), .Q(n5084), .QN(net86699) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n2776), .CK(CLK), .QN(n4024) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n2775), .CK(CLK), .QN(n4042) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n2774), .CK(CLK), .QN(n4060) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n2773), .CK(CLK), .QN(n4078) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n2772), .CK(CLK), .QN(n4114) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n2771), .CK(CLK), .QN(n4132) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n2770), .CK(CLK), .QN(n4150) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n2769), .CK(CLK), .QN(n4168) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n2768), .CK(CLK), .QN(n4186) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n2767), .CK(CLK), .QN(n4204) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n2766), .CK(CLK), .QN(n4222) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n2765), .CK(CLK), .QN(n4240) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n2764), .CK(CLK), .QN(n4258) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n2763), .CK(CLK), .QN(n4276) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n2762), .CK(CLK), .QN(n3736) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n2761), .CK(CLK), .QN(n3754) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n2760), .CK(CLK), .QN(n3772) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n2759), .CK(CLK), .QN(n3790) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n2758), .CK(CLK), .QN(n3808) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n2757), .CK(CLK), .QN(n3826) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n2756), .CK(CLK), .QN(n3844) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n2755), .CK(CLK), .QN(n3898) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n2754), .CK(CLK), .QN(n4096) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n2753), .CK(CLK), .QN(n4294) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n2744), .CK(CLK), .QN(n4025) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n2743), .CK(CLK), .QN(n4043) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n2742), .CK(CLK), .QN(n4061) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n2741), .CK(CLK), .QN(n4079) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n2740), .CK(CLK), .QN(n4115) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n2739), .CK(CLK), .QN(n4133) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n2738), .CK(CLK), .QN(n4151) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n2737), .CK(CLK), .QN(n4169) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n2736), .CK(CLK), .QN(n4187) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n2735), .CK(CLK), .QN(n4205) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n2734), .CK(CLK), .QN(n4223) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n2733), .CK(CLK), .QN(n4241) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n2732), .CK(CLK), .QN(n4259) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n2731), .CK(CLK), .QN(n4277) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n2730), .CK(CLK), .QN(n3737) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n2729), .CK(CLK), .QN(n3755) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n2728), .CK(CLK), .QN(n3773) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n2727), .CK(CLK), .QN(n3791) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n2726), .CK(CLK), .QN(n3809) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n2725), .CK(CLK), .QN(n3827) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n2724), .CK(CLK), .QN(n3845) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n2723), .CK(CLK), .QN(n3899) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n2722), .CK(CLK), .QN(n4097) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n2721), .CK(CLK), .QN(n4295) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n3660), .CK(CLK), .QN(n428) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n3659), .CK(CLK), .QN(n435) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n3649), .CK(CLK), .QN(n442) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n2808), .CK(CLK), .Q(n4554), .QN(
        net86754) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2807), .CK(CLK), .Q(n4588), .QN(
        net86753) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n2806), .CK(CLK), .Q(n4622), .QN(
        net86752) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2805), .CK(CLK), .Q(n4656), .QN(
        net86751) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n2804), .CK(CLK), .Q(n4724), .QN(
        net86750) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n2803), .CK(CLK), .Q(n4758), .QN(
        net86749) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n2802), .CK(CLK), .Q(n4792), .QN(
        net86748) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n2801), .CK(CLK), .Q(n4826), .QN(
        net86747) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n2800), .CK(CLK), .Q(n4860), .QN(
        net86746) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n2799), .CK(CLK), .Q(n4894), .QN(
        net86745) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n2798), .CK(CLK), .Q(n4928), .QN(
        net86744) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n2797), .CK(CLK), .Q(n4962), .QN(
        net86743) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n2796), .CK(CLK), .Q(n4996), .QN(
        net86742) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2795), .CK(CLK), .Q(n5030), .QN(
        net86741) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n2794), .CK(CLK), .Q(n2404), .QN(net86740) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n2793), .CK(CLK), .Q(n2443), .QN(net86739) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n2792), .CK(CLK), .Q(n2477), .QN(net86738) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2791), .CK(CLK), .Q(n2511), .QN(net86737) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2790), .CK(CLK), .Q(n2545), .QN(net86736) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n2789), .CK(CLK), .Q(n2579), .QN(net86735) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2788), .CK(CLK), .Q(n2613), .QN(net86734) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n2787), .CK(CLK), .Q(n4316), .QN(net86733) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n2786), .CK(CLK), .Q(n4690), .QN(net86732) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n2785), .CK(CLK), .Q(n5077), .QN(net86731) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n2840), .CK(CLK), .Q(n4555), .QN(
        net86786) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n2839), .CK(CLK), .Q(n4589), .QN(
        net86785) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n2838), .CK(CLK), .Q(n4623), .QN(
        net86784) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n2837), .CK(CLK), .Q(n4657), .QN(
        net86783) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n2836), .CK(CLK), .Q(n4725), .QN(
        net86782) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n2835), .CK(CLK), .Q(n4759), .QN(
        net86781) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n2834), .CK(CLK), .Q(n4793), .QN(
        net86780) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n2833), .CK(CLK), .Q(n4827), .QN(
        net86779) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n2832), .CK(CLK), .Q(n4861), .QN(
        net86778) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n2831), .CK(CLK), .Q(n4895), .QN(
        net86777) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n2830), .CK(CLK), .Q(n4929), .QN(
        net86776) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n2829), .CK(CLK), .Q(n4963), .QN(
        net86775) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n2828), .CK(CLK), .Q(n4997), .QN(
        net86774) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2827), .CK(CLK), .Q(n5031), .QN(
        net86773) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n2826), .CK(CLK), .Q(n2406), .QN(net86772) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n2825), .CK(CLK), .Q(n2444), .QN(net86771) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n2824), .CK(CLK), .Q(n2478), .QN(net86770) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2823), .CK(CLK), .Q(n2512), .QN(net86769) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2822), .CK(CLK), .Q(n2546), .QN(net86768) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n2821), .CK(CLK), .Q(n2580), .QN(net86767) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2820), .CK(CLK), .Q(n2614), .QN(net86766) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n2819), .CK(CLK), .Q(n4317), .QN(net86765) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n2818), .CK(CLK), .Q(n4691), .QN(net86764) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n2817), .CK(CLK), .Q(n5078), .QN(net86763) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n2936), .CK(CLK), .Q(n4548), .QN(
        net86818) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n2935), .CK(CLK), .Q(n4582), .QN(
        net86817) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n2934), .CK(CLK), .Q(n4616), .QN(
        net86816) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n2933), .CK(CLK), .Q(n4650), .QN(
        net86815) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n2932), .CK(CLK), .Q(n4718), .QN(
        net86814) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n2931), .CK(CLK), .Q(n4752), .QN(
        net86813) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n2930), .CK(CLK), .Q(n4786), .QN(
        net86812) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n2929), .CK(CLK), .Q(n4820), .QN(
        net86811) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n2928), .CK(CLK), .Q(n4854), .QN(
        net86810) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n2927), .CK(CLK), .Q(n4888), .QN(
        net86809) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n2926), .CK(CLK), .Q(n4922), .QN(
        net86808) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n2925), .CK(CLK), .Q(n4956), .QN(
        net86807) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n2924), .CK(CLK), .Q(n4990), .QN(
        net86806) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n2923), .CK(CLK), .Q(n5024), .QN(
        net86805) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n2922), .CK(CLK), .Q(n2390), .QN(net86804) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n2921), .CK(CLK), .Q(n2437), .QN(net86803) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n2920), .CK(CLK), .Q(n2471), .QN(net86802) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n2919), .CK(CLK), .Q(n2505), .QN(net86801) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n2918), .CK(CLK), .Q(n2539), .QN(net86800) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n2917), .CK(CLK), .Q(n2573), .QN(net86799) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n2916), .CK(CLK), .Q(n2607), .QN(net86798) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n2915), .CK(CLK), .Q(n4310), .QN(net86797) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n2914), .CK(CLK), .Q(n4684), .QN(net86796) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n2913), .CK(CLK), .Q(n5068), .QN(net86795) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n2968), .CK(CLK), .Q(n4549), .QN(
        net86850) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n2967), .CK(CLK), .Q(n4583), .QN(
        net86849) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n2966), .CK(CLK), .Q(n4617), .QN(
        net86848) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n2965), .CK(CLK), .Q(n4651), .QN(
        net86847) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n2964), .CK(CLK), .Q(n4719), .QN(
        net86846) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n2963), .CK(CLK), .Q(n4753), .QN(
        net86845) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n2962), .CK(CLK), .Q(n4787), .QN(
        net86844) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n2961), .CK(CLK), .Q(n4821), .QN(
        net86843) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n2960), .CK(CLK), .Q(n4855), .QN(
        net86842) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n2959), .CK(CLK), .Q(n4889), .QN(
        net86841) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n2958), .CK(CLK), .Q(n4923), .QN(
        net86840) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n2957), .CK(CLK), .Q(n4957), .QN(
        net86839) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n2956), .CK(CLK), .Q(n4991), .QN(
        net86838) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n2955), .CK(CLK), .Q(n5025), .QN(
        net86837) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n2954), .CK(CLK), .Q(n2392), .QN(net86836) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n2953), .CK(CLK), .Q(n2438), .QN(net86835) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n2952), .CK(CLK), .Q(n2472), .QN(net86834) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n2951), .CK(CLK), .Q(n2506), .QN(net86833) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n2950), .CK(CLK), .Q(n2540), .QN(net86832) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n2949), .CK(CLK), .Q(n2574), .QN(net86831) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n2948), .CK(CLK), .Q(n2608), .QN(net86830) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n2947), .CK(CLK), .Q(n4311), .QN(net86829) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n2946), .CK(CLK), .Q(n4685), .QN(net86828) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n2945), .CK(CLK), .Q(n5069), .QN(net86827) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n3064), .CK(CLK), .Q(n4551), .QN(
        net86882) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n3063), .CK(CLK), .Q(n4585), .QN(
        net86881) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n3062), .CK(CLK), .Q(n4619), .QN(
        net86880) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n3061), .CK(CLK), .Q(n4653), .QN(
        net86879) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n3060), .CK(CLK), .Q(n4721), .QN(
        net86878) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n3059), .CK(CLK), .Q(n4755), .QN(
        net86877) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n3058), .CK(CLK), .Q(n4789), .QN(
        net86876) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n3057), .CK(CLK), .Q(n4823), .QN(
        net86875) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n3056), .CK(CLK), .Q(n4857), .QN(
        net86874) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n3055), .CK(CLK), .Q(n4891), .QN(
        net86873) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n3054), .CK(CLK), .Q(n4925), .QN(
        net86872) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n3053), .CK(CLK), .Q(n4959), .QN(
        net86871) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n3052), .CK(CLK), .Q(n4993), .QN(
        net86870) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n3051), .CK(CLK), .Q(n5027), .QN(
        net86869) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n3050), .CK(CLK), .Q(n2397), .QN(net86868) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n3049), .CK(CLK), .Q(n2440), .QN(net86867) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n3048), .CK(CLK), .Q(n2474), .QN(net86866) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n3047), .CK(CLK), .Q(n2508), .QN(net86865) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n3046), .CK(CLK), .Q(n2542), .QN(net86864) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n3045), .CK(CLK), .Q(n2576), .QN(net86863) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n3044), .CK(CLK), .Q(n2610), .QN(net86862) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n3043), .CK(CLK), .Q(n4313), .QN(net86861) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n3042), .CK(CLK), .Q(n4687), .QN(net86860) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n3041), .CK(CLK), .Q(n5073), .QN(net86859) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n3096), .CK(CLK), .Q(n4552), .QN(
        net86914) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n3095), .CK(CLK), .Q(n4586), .QN(
        net86913) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n3094), .CK(CLK), .Q(n4620), .QN(
        net86912) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n3093), .CK(CLK), .Q(n4654), .QN(
        net86911) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n3092), .CK(CLK), .Q(n4722), .QN(
        net86910) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n3091), .CK(CLK), .Q(n4756), .QN(
        net86909) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n3090), .CK(CLK), .Q(n4790), .QN(
        net86908) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n3089), .CK(CLK), .Q(n4824), .QN(
        net86907) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n3088), .CK(CLK), .Q(n4858), .QN(
        net86906) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n3087), .CK(CLK), .Q(n4892), .QN(
        net86905) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n3086), .CK(CLK), .Q(n4926), .QN(
        net86904) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n3085), .CK(CLK), .Q(n4960), .QN(
        net86903) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n3084), .CK(CLK), .Q(n4994), .QN(
        net86902) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n3083), .CK(CLK), .Q(n5028), .QN(
        net86901) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n3082), .CK(CLK), .Q(n2399), .QN(net86900) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n3081), .CK(CLK), .Q(n2441), .QN(net86899) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n3080), .CK(CLK), .Q(n2475), .QN(net86898) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n3079), .CK(CLK), .Q(n2509), .QN(net86897) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n3078), .CK(CLK), .Q(n2543), .QN(net86896) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n3077), .CK(CLK), .Q(n2577), .QN(net86895) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n3076), .CK(CLK), .Q(n2611), .QN(net86894) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n3075), .CK(CLK), .Q(n4314), .QN(net86893) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n3074), .CK(CLK), .Q(n4688), .QN(net86892) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n3073), .CK(CLK), .Q(n5074), .QN(net86891) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n3192), .CK(CLK), .Q(n4533), .QN(
        net86946) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n3191), .CK(CLK), .Q(n4567), .QN(
        net86945) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n3190), .CK(CLK), .Q(n4601), .QN(
        net86944) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n3189), .CK(CLK), .Q(n4635), .QN(
        net86943) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n3188), .CK(CLK), .Q(n4703), .QN(
        net86942) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n3187), .CK(CLK), .Q(n4737), .QN(
        net86941) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n3186), .CK(CLK), .Q(n4771), .QN(
        net86940) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n3185), .CK(CLK), .Q(n4805), .QN(
        net86939) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n3184), .CK(CLK), .Q(n4839), .QN(
        net86938) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n3183), .CK(CLK), .Q(n4873), .QN(
        net86937) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n3182), .CK(CLK), .Q(n4907), .QN(
        net86936) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n3181), .CK(CLK), .Q(n4941), .QN(
        net86935) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n3180), .CK(CLK), .Q(n4975), .QN(
        net86934) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n3179), .CK(CLK), .Q(n5009), .QN(
        net86933) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n3178), .CK(CLK), .Q(n2360), .QN(net86932) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n3177), .CK(CLK), .Q(n2422), .QN(net86931) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n3176), .CK(CLK), .Q(n2456), .QN(net86930) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n3175), .CK(CLK), .Q(n2490), .QN(net86929) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n3174), .CK(CLK), .Q(n2524), .QN(net86928) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n3173), .CK(CLK), .Q(n2558), .QN(net86927) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n3172), .CK(CLK), .Q(n2592), .QN(net86926) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n3171), .CK(CLK), .Q(n3719), .QN(net86925) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n3170), .CK(CLK), .Q(n4669), .QN(net86924) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n3169), .CK(CLK), .Q(n5043), .QN(net86923) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n3224), .CK(CLK), .Q(n4532), .QN(
        net86978) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n3223), .CK(CLK), .Q(n4566), .QN(
        net86977) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n3222), .CK(CLK), .Q(n4600), .QN(
        net86976) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n3221), .CK(CLK), .Q(n4634), .QN(
        net86975) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n3220), .CK(CLK), .Q(n4702), .QN(
        net86974) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n3219), .CK(CLK), .Q(n4736), .QN(
        net86973) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n3218), .CK(CLK), .Q(n4770), .QN(
        net86972) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n3217), .CK(CLK), .Q(n4804), .QN(
        net86971) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n3216), .CK(CLK), .Q(n4838), .QN(
        net86970) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n3215), .CK(CLK), .Q(n4872), .QN(
        net86969) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n3214), .CK(CLK), .Q(n4906), .QN(
        net86968) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n3213), .CK(CLK), .Q(n4940), .QN(
        net86967) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n3212), .CK(CLK), .Q(n4974), .QN(
        net86966) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n3211), .CK(CLK), .Q(n5008), .QN(
        net86965) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n3210), .CK(CLK), .Q(n2358), .QN(net86964) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n3209), .CK(CLK), .Q(n2421), .QN(net86963) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n3208), .CK(CLK), .Q(n2455), .QN(net86962) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n3207), .CK(CLK), .Q(n2489), .QN(net86961) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n3206), .CK(CLK), .Q(n2523), .QN(net86960) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n3205), .CK(CLK), .Q(n2557), .QN(net86959) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n3204), .CK(CLK), .Q(n2591), .QN(net86958) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n3203), .CK(CLK), .Q(n3718), .QN(net86957) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n3202), .CK(CLK), .Q(n4668), .QN(net86956) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n3201), .CK(CLK), .Q(n5042), .QN(net86955) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n3320), .CK(CLK), .Q(n4536), .QN(
        net87010) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n3319), .CK(CLK), .Q(n4570), .QN(
        net87009) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n3318), .CK(CLK), .Q(n4604), .QN(
        net87008) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n3317), .CK(CLK), .Q(n4638), .QN(
        net87007) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n3316), .CK(CLK), .Q(n4706), .QN(
        net87006) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n3315), .CK(CLK), .Q(n4740), .QN(
        net87005) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n3314), .CK(CLK), .Q(n4774), .QN(
        net87004) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n3313), .CK(CLK), .Q(n4808), .QN(
        net87003) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n3312), .CK(CLK), .Q(n4842), .QN(
        net87002) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n3311), .CK(CLK), .Q(n4876), .QN(
        net87001) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n3310), .CK(CLK), .Q(n4910), .QN(
        net87000) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n3309), .CK(CLK), .Q(n4944), .QN(
        net86999) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n3308), .CK(CLK), .Q(n4978), .QN(
        net86998) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n3307), .CK(CLK), .Q(n5012), .QN(
        net86997) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n3306), .CK(CLK), .Q(n2367), .QN(net86996) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n3305), .CK(CLK), .Q(n2425), .QN(net86995) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n3304), .CK(CLK), .Q(n2459), .QN(net86994) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n3303), .CK(CLK), .Q(n2493), .QN(net86993) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n3302), .CK(CLK), .Q(n2527), .QN(net86992) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n3301), .CK(CLK), .Q(n2561), .QN(net86991) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n3300), .CK(CLK), .Q(n2595), .QN(net86990) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n3299), .CK(CLK), .Q(n4298), .QN(net86989) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n3298), .CK(CLK), .Q(n4672), .QN(net86988) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n3297), .CK(CLK), .Q(n5050), .QN(net86987) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n3352), .CK(CLK), .Q(n4535), .QN(
        net87042) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n3351), .CK(CLK), .Q(n4569), .QN(
        net87041) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n3350), .CK(CLK), .Q(n4603), .QN(
        net87040) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n3349), .CK(CLK), .Q(n4637), .QN(
        net87039) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n3348), .CK(CLK), .Q(n4705), .QN(
        net87038) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n3347), .CK(CLK), .Q(n4739), .QN(
        net87037) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n3346), .CK(CLK), .Q(n4773), .QN(
        net87036) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n3345), .CK(CLK), .Q(n4807), .QN(
        net87035) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n3344), .CK(CLK), .Q(n4841), .QN(
        net87034) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n3343), .CK(CLK), .Q(n4875), .QN(
        net87033) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n3342), .CK(CLK), .Q(n4909), .QN(
        net87032) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n3341), .CK(CLK), .Q(n4943), .QN(
        net87031) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n3340), .CK(CLK), .Q(n4977), .QN(
        net87030) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n3339), .CK(CLK), .Q(n5011), .QN(
        net87029) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n3338), .CK(CLK), .Q(n2365), .QN(net87028) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n3337), .CK(CLK), .Q(n2424), .QN(net87027) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n3336), .CK(CLK), .Q(n2458), .QN(net87026) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n3335), .CK(CLK), .Q(n2492), .QN(net87025) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n3334), .CK(CLK), .Q(n2526), .QN(net87024) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n3333), .CK(CLK), .Q(n2560), .QN(net87023) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n3332), .CK(CLK), .Q(n2594), .QN(net87022) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n3331), .CK(CLK), .Q(n3721), .QN(net87021) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n3330), .CK(CLK), .Q(n4671), .QN(net87020) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n3329), .CK(CLK), .Q(n5049), .QN(net87019) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n3448), .CK(CLK), .Q(n4539), .QN(net87074) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n3447), .CK(CLK), .Q(n4573), .QN(net87073) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n3446), .CK(CLK), .Q(n4607), .QN(net87072) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n3445), .CK(CLK), .Q(n4641), .QN(net87071) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n3444), .CK(CLK), .Q(n4709), .QN(net87070) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n3443), .CK(CLK), .Q(n4743), .QN(net87069) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n3442), .CK(CLK), .Q(n4777), .QN(net87068) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n3441), .CK(CLK), .Q(n4811), .QN(net87067) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n3440), .CK(CLK), .Q(n4845), .QN(net87066) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n3439), .CK(CLK), .Q(n4879), .QN(net87065) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n3438), .CK(CLK), .Q(n4913), .QN(net87064) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n3437), .CK(CLK), .Q(n4947), .QN(net87063) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n3436), .CK(CLK), .Q(n4981), .QN(net87062) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n3435), .CK(CLK), .Q(n5015), .QN(net87061) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n3434), .CK(CLK), .Q(n2374), .QN(net87060)
         );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n3433), .CK(CLK), .Q(n2428), .QN(net87059)
         );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n3432), .CK(CLK), .Q(n2462), .QN(net87058)
         );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n3431), .CK(CLK), .Q(n2496), .QN(net87057)
         );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n3430), .CK(CLK), .Q(n2530), .QN(net87056)
         );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n3429), .CK(CLK), .Q(n2564), .QN(net87055)
         );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n3428), .CK(CLK), .Q(n2598), .QN(net87054)
         );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n3427), .CK(CLK), .Q(n4301), .QN(net87053)
         );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n3426), .CK(CLK), .Q(n4675), .QN(net87052)
         );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n3425), .CK(CLK), .Q(n5057), .QN(net87051)
         );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n3480), .CK(CLK), .Q(n4538), .QN(net87106) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n3479), .CK(CLK), .Q(n4572), .QN(net87105) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n3478), .CK(CLK), .Q(n4606), .QN(net87104) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n3477), .CK(CLK), .Q(n4640), .QN(net87103) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n3476), .CK(CLK), .Q(n4708), .QN(net87102) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n3475), .CK(CLK), .Q(n4742), .QN(net87101) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n3474), .CK(CLK), .Q(n4776), .QN(net87100) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n3473), .CK(CLK), .Q(n4810), .QN(net87099) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n3472), .CK(CLK), .Q(n4844), .QN(net87098) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n3471), .CK(CLK), .Q(n4878), .QN(net87097) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n3470), .CK(CLK), .Q(n4912), .QN(net87096) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n3469), .CK(CLK), .Q(n4946), .QN(net87095) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n3468), .CK(CLK), .Q(n4980), .QN(net87094) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n3467), .CK(CLK), .Q(n5014), .QN(net87093) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n3466), .CK(CLK), .Q(n2372), .QN(net87092)
         );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n3465), .CK(CLK), .Q(n2427), .QN(net87091)
         );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n3464), .CK(CLK), .Q(n2461), .QN(net87090)
         );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n3463), .CK(CLK), .Q(n2495), .QN(net87089)
         );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n3462), .CK(CLK), .Q(n2529), .QN(net87088)
         );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n3461), .CK(CLK), .Q(n2563), .QN(net87087)
         );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n3460), .CK(CLK), .Q(n2597), .QN(net87086)
         );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n3459), .CK(CLK), .Q(n4300), .QN(net87085)
         );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n3458), .CK(CLK), .Q(n4674), .QN(net87084)
         );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n3457), .CK(CLK), .Q(n5056), .QN(net87083)
         );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n2880), .CK(CLK), .QN(n54) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n2879), .CK(CLK), .QN(n61) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n2878), .CK(CLK), .QN(n75) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n2877), .CK(CLK), .QN(n82) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n2876), .CK(CLK), .QN(n89) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n2875), .CK(CLK), .QN(n96) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n2858), .CK(CLK), .QN(n5) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n2853), .CK(CLK), .QN(n40) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n2852), .CK(CLK), .QN(n47) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n2851), .CK(CLK), .QN(n68) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n3040), .CK(CLK), .QN(n56) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n3039), .CK(CLK), .QN(n63) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n3038), .CK(CLK), .QN(n77) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n3037), .CK(CLK), .QN(n84) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n3036), .CK(CLK), .QN(n91) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n3035), .CK(CLK), .QN(n98) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n3018), .CK(CLK), .QN(n7) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n3013), .CK(CLK), .QN(n42) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n3012), .CK(CLK), .QN(n49) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n3011), .CK(CLK), .QN(n70) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n3168), .CK(CLK), .QN(n55) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n3167), .CK(CLK), .QN(n62) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n3166), .CK(CLK), .QN(n76) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n3165), .CK(CLK), .QN(n83) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n3164), .CK(CLK), .QN(n90) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n3163), .CK(CLK), .QN(n97) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n3146), .CK(CLK), .QN(n6) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n3141), .CK(CLK), .QN(n41) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n3140), .CK(CLK), .QN(n48) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n3139), .CK(CLK), .QN(n69) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n3264), .CK(CLK), .QN(n53) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n3263), .CK(CLK), .QN(n60) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n3262), .CK(CLK), .QN(n74) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n3261), .CK(CLK), .QN(n81) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n3260), .CK(CLK), .QN(n88) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n3259), .CK(CLK), .QN(n95) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n3242), .CK(CLK), .QN(n4) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n3237), .CK(CLK), .QN(n39) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n3236), .CK(CLK), .QN(n46) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n3235), .CK(CLK), .QN(n67) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n3520), .CK(CLK), .QN(n51) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n3519), .CK(CLK), .QN(n58) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n3518), .CK(CLK), .QN(n72) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n3517), .CK(CLK), .QN(n79) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n3516), .CK(CLK), .QN(n86) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n3515), .CK(CLK), .QN(n93) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n3497), .CK(CLK), .QN(n9) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n3492), .CK(CLK), .QN(n44) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n3491), .CK(CLK), .QN(n65) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n3392), .CK(CLK), .QN(n52) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n3391), .CK(CLK), .QN(n59) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n3390), .CK(CLK), .QN(n73) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n3389), .CK(CLK), .QN(n80) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n3388), .CK(CLK), .QN(n87) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n3387), .CK(CLK), .QN(n94) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n3364), .CK(CLK), .QN(n45) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n3363), .CK(CLK), .QN(n66) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n3608), .CK(CLK), .Q(n4541), .QN(net87170) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n3607), .CK(CLK), .Q(n4575), .QN(net87169) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n3606), .CK(CLK), .Q(n4609), .QN(net87168) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n3605), .CK(CLK), .Q(n4643), .QN(net87167) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n3604), .CK(CLK), .Q(n4711), .QN(net87166) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n3603), .CK(CLK), .Q(n4745), .QN(net87165) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n3602), .CK(CLK), .Q(n4779), .QN(net87164) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n3601), .CK(CLK), .Q(n4813), .QN(net87163) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n3600), .CK(CLK), .Q(n4847), .QN(net87162) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n3599), .CK(CLK), .Q(n4881), .QN(net87161) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n3598), .CK(CLK), .Q(n4915), .QN(net87160) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n3597), .CK(CLK), .Q(n4949), .QN(net87159) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n3596), .CK(CLK), .Q(n4983), .QN(net87158) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n3595), .CK(CLK), .Q(n5017), .QN(net87157) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n3594), .CK(CLK), .Q(n2379), .QN(net87156)
         );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n3593), .CK(CLK), .Q(n2430), .QN(net87155)
         );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n3592), .CK(CLK), .Q(n2464), .QN(net87154)
         );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n3591), .CK(CLK), .Q(n2498), .QN(net87153)
         );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n3590), .CK(CLK), .Q(n2532), .QN(net87152)
         );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n3589), .CK(CLK), .Q(n2566), .QN(net87151)
         );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n3588), .CK(CLK), .Q(n2600), .QN(net87150)
         );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n3587), .CK(CLK), .Q(n4303), .QN(net87149)
         );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n3586), .CK(CLK), .Q(n4677), .QN(net87148)
         );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n3585), .CK(CLK), .Q(n5061), .QN(net87147)
         );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n3576), .CK(CLK), .Q(n4542), .QN(net87138) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n3575), .CK(CLK), .Q(n4576), .QN(net87137) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n3574), .CK(CLK), .Q(n4610), .QN(net87136) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n3573), .CK(CLK), .Q(n4644), .QN(net87135) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n3572), .CK(CLK), .Q(n4712), .QN(net87134) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n3571), .CK(CLK), .Q(n4746), .QN(net87133) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n3570), .CK(CLK), .Q(n4780), .QN(net87132) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n3569), .CK(CLK), .Q(n4814), .QN(net87131) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n3568), .CK(CLK), .Q(n4848), .QN(net87130) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n3567), .CK(CLK), .Q(n4882), .QN(net87129) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n3566), .CK(CLK), .Q(n4916), .QN(net87128) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n3565), .CK(CLK), .Q(n4950), .QN(net87127) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n3564), .CK(CLK), .Q(n4984), .QN(net87126) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n3563), .CK(CLK), .Q(n5018), .QN(net87125) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n3562), .CK(CLK), .Q(n2381), .QN(net87124)
         );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n3561), .CK(CLK), .Q(n2431), .QN(net87123)
         );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n3560), .CK(CLK), .Q(n2465), .QN(net87122)
         );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n3559), .CK(CLK), .Q(n2499), .QN(net87121)
         );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n3558), .CK(CLK), .Q(n2533), .QN(net87120)
         );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n3557), .CK(CLK), .Q(n2567), .QN(net87119)
         );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n3556), .CK(CLK), .Q(n2601), .QN(net87118)
         );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n3555), .CK(CLK), .Q(n4304), .QN(net87117)
         );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n3554), .CK(CLK), .Q(n4678), .QN(net87116)
         );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n3553), .CK(CLK), .Q(n5062), .QN(net87115)
         );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n2893), .CK(CLK), .QN(n425) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n2892), .CK(CLK), .QN(n432) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n2891), .CK(CLK), .QN(n439) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n2881), .CK(CLK), .QN(n446) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n2989), .CK(CLK), .QN(n427) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n2988), .CK(CLK), .QN(n434) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n2987), .CK(CLK), .QN(n441) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n2977), .CK(CLK), .QN(n448) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n3117), .CK(CLK), .QN(n426) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n3116), .CK(CLK), .QN(n433) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n3115), .CK(CLK), .QN(n440) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n3105), .CK(CLK), .QN(n447) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n3277), .CK(CLK), .QN(n424) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n3276), .CK(CLK), .QN(n431) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n3275), .CK(CLK), .QN(n438) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n3265), .CK(CLK), .QN(n445) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n3405), .CK(CLK), .QN(n423) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n3404), .CK(CLK), .QN(n430) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n3403), .CK(CLK), .QN(n437) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n3393), .CK(CLK), .QN(n444) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n3532), .CK(CLK), .QN(n429) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n3531), .CK(CLK), .QN(n436) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n3521), .CK(CLK), .QN(n443) );
  NOR3_X1 U3 ( .A1(n5691), .A2(ADD_RD1[4]), .A3(n5692), .ZN(n5684) );
  NOR3_X1 U4 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n5692), .ZN(n5686) );
  NOR3_X1 U5 ( .A1(n5053), .A2(ADD_RD2[4]), .A3(n5054), .ZN(n5044) );
  NOR3_X1 U6 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n5054), .ZN(n5046) );
  INV_X1 U7 ( .A(n6492), .ZN(n6485) );
  INV_X1 U8 ( .A(n6729), .ZN(n6722) );
  INV_X1 U9 ( .A(n6357), .ZN(n6348) );
  INV_X1 U10 ( .A(n6411), .ZN(n6404) );
  INV_X1 U11 ( .A(n6420), .ZN(n6413) );
  INV_X1 U12 ( .A(n6447), .ZN(n6440) );
  INV_X1 U13 ( .A(n6456), .ZN(n6449) );
  INV_X1 U14 ( .A(n6483), .ZN(n6476) );
  INV_X1 U15 ( .A(n6519), .ZN(n6512) );
  INV_X1 U16 ( .A(n6528), .ZN(n6521) );
  INV_X1 U17 ( .A(n6555), .ZN(n6548) );
  INV_X1 U18 ( .A(n6564), .ZN(n6557) );
  INV_X1 U19 ( .A(n6591), .ZN(n6584) );
  INV_X1 U20 ( .A(n6600), .ZN(n6593) );
  INV_X1 U21 ( .A(n6627), .ZN(n6620) );
  INV_X1 U22 ( .A(n6366), .ZN(n6359) );
  INV_X1 U23 ( .A(n6375), .ZN(n6368) );
  INV_X1 U24 ( .A(n6384), .ZN(n6377) );
  INV_X1 U25 ( .A(n6393), .ZN(n6386) );
  INV_X1 U26 ( .A(n6402), .ZN(n6395) );
  INV_X1 U27 ( .A(n6429), .ZN(n6422) );
  INV_X1 U28 ( .A(n6438), .ZN(n6431) );
  INV_X1 U29 ( .A(n6465), .ZN(n6458) );
  INV_X1 U30 ( .A(n6474), .ZN(n6467) );
  INV_X1 U31 ( .A(n6501), .ZN(n6494) );
  INV_X1 U32 ( .A(n6510), .ZN(n6503) );
  INV_X1 U33 ( .A(n6537), .ZN(n6530) );
  INV_X1 U34 ( .A(n6546), .ZN(n6539) );
  INV_X1 U35 ( .A(n6573), .ZN(n6566) );
  INV_X1 U36 ( .A(n6582), .ZN(n6575) );
  INV_X1 U37 ( .A(n6609), .ZN(n6602) );
  INV_X1 U38 ( .A(n6618), .ZN(n6611) );
  INV_X1 U39 ( .A(RESET), .ZN(n6736) );
  BUF_X1 U40 ( .A(n6493), .Z(n6486) );
  BUF_X1 U41 ( .A(n6493), .Z(n6487) );
  BUF_X1 U42 ( .A(n6493), .Z(n6488) );
  BUF_X1 U43 ( .A(n6493), .Z(n6489) );
  BUF_X1 U44 ( .A(n6493), .Z(n6490) );
  BUF_X1 U45 ( .A(n6493), .Z(n6491) );
  BUF_X1 U46 ( .A(n6730), .Z(n6723) );
  BUF_X1 U47 ( .A(n6730), .Z(n6724) );
  BUF_X1 U48 ( .A(n6730), .Z(n6725) );
  BUF_X1 U49 ( .A(n6730), .Z(n6726) );
  BUF_X1 U50 ( .A(n6730), .Z(n6727) );
  BUF_X1 U51 ( .A(n6730), .Z(n6728) );
  BUF_X1 U52 ( .A(n6493), .Z(n6492) );
  BUF_X1 U53 ( .A(n6730), .Z(n6729) );
  BUF_X1 U54 ( .A(n6358), .Z(n6357) );
  BUF_X1 U55 ( .A(n6351), .Z(n6355) );
  BUF_X1 U56 ( .A(n6358), .Z(n6354) );
  BUF_X1 U57 ( .A(n6358), .Z(n6353) );
  BUF_X1 U58 ( .A(n6358), .Z(n6352) );
  BUF_X1 U59 ( .A(n6358), .Z(n6351) );
  BUF_X1 U60 ( .A(n6358), .Z(n6350) );
  BUF_X1 U61 ( .A(n6358), .Z(n6349) );
  BUF_X1 U62 ( .A(n6350), .Z(n6356) );
  INV_X1 U63 ( .A(n5103), .ZN(n6044) );
  INV_X1 U64 ( .A(n5104), .ZN(n6052) );
  INV_X1 U65 ( .A(n5108), .ZN(n6012) );
  INV_X1 U66 ( .A(n5109), .ZN(n6020) );
  INV_X1 U67 ( .A(n5108), .ZN(n6013) );
  AND2_X1 U68 ( .A1(n5708), .A2(n5685), .ZN(n5136) );
  INV_X1 U69 ( .A(n5093), .ZN(n6096) );
  INV_X1 U70 ( .A(n5098), .ZN(n6076) );
  INV_X1 U71 ( .A(n5099), .ZN(n6084) );
  INV_X1 U72 ( .A(n5094), .ZN(n6104) );
  INV_X1 U73 ( .A(n5098), .ZN(n6077) );
  INV_X1 U74 ( .A(n5094), .ZN(n6105) );
  INV_X1 U75 ( .A(n5099), .ZN(n6085) );
  INV_X1 U76 ( .A(n5127), .ZN(n5916) );
  INV_X1 U77 ( .A(n5133), .ZN(n5892) );
  INV_X1 U78 ( .A(n5117), .ZN(n5980) );
  INV_X1 U79 ( .A(n5118), .ZN(n5988) );
  INV_X1 U80 ( .A(n5122), .ZN(n5948) );
  INV_X1 U81 ( .A(n5123), .ZN(n5956) );
  INV_X1 U82 ( .A(n5127), .ZN(n5917) );
  INV_X1 U83 ( .A(n5128), .ZN(n5924) );
  INV_X1 U84 ( .A(n5133), .ZN(n5893) );
  INV_X1 U85 ( .A(n5118), .ZN(n5989) );
  INV_X1 U86 ( .A(n5123), .ZN(n5957) );
  INV_X1 U87 ( .A(n5132), .ZN(n5884) );
  INV_X1 U88 ( .A(n5117), .ZN(n5981) );
  INV_X1 U89 ( .A(n5122), .ZN(n5949) );
  INV_X1 U90 ( .A(n1880), .ZN(n6730) );
  OAI21_X1 U91 ( .B1(n1941), .B2(n1942), .A(n6735), .ZN(n1880) );
  BUF_X1 U92 ( .A(n1902), .Z(n6690) );
  BUF_X1 U93 ( .A(n1900), .Z(n6693) );
  BUF_X1 U94 ( .A(n1898), .Z(n6696) );
  BUF_X1 U95 ( .A(n1896), .Z(n6699) );
  BUF_X1 U96 ( .A(n1894), .Z(n6702) );
  BUF_X1 U97 ( .A(n1892), .Z(n6705) );
  BUF_X1 U98 ( .A(n1890), .Z(n6708) );
  BUF_X1 U99 ( .A(n1888), .Z(n6711) );
  BUF_X1 U100 ( .A(n1886), .Z(n6714) );
  BUF_X1 U101 ( .A(n1884), .Z(n6717) );
  BUF_X1 U102 ( .A(n1882), .Z(n6720) );
  BUF_X1 U103 ( .A(n1879), .Z(n6732) );
  BUF_X1 U104 ( .A(n1902), .Z(n6689) );
  BUF_X1 U105 ( .A(n1900), .Z(n6692) );
  BUF_X1 U106 ( .A(n1898), .Z(n6695) );
  BUF_X1 U107 ( .A(n1896), .Z(n6698) );
  BUF_X1 U108 ( .A(n1894), .Z(n6701) );
  BUF_X1 U109 ( .A(n1892), .Z(n6704) );
  BUF_X1 U110 ( .A(n1890), .Z(n6707) );
  BUF_X1 U111 ( .A(n1888), .Z(n6710) );
  BUF_X1 U112 ( .A(n1886), .Z(n6713) );
  BUF_X1 U113 ( .A(n1884), .Z(n6716) );
  BUF_X1 U114 ( .A(n1882), .Z(n6719) );
  BUF_X1 U115 ( .A(n1879), .Z(n6731) );
  BUF_X1 U116 ( .A(n1940), .Z(n6629) );
  BUF_X1 U117 ( .A(n1938), .Z(n6633) );
  BUF_X1 U118 ( .A(n1936), .Z(n6636) );
  BUF_X1 U119 ( .A(n1934), .Z(n6639) );
  BUF_X1 U120 ( .A(n1932), .Z(n6642) );
  BUF_X1 U121 ( .A(n1930), .Z(n6645) );
  BUF_X1 U122 ( .A(n1928), .Z(n6648) );
  BUF_X1 U123 ( .A(n1926), .Z(n6651) );
  BUF_X1 U124 ( .A(n1924), .Z(n6654) );
  BUF_X1 U125 ( .A(n1922), .Z(n6657) );
  BUF_X1 U126 ( .A(n1921), .Z(n6660) );
  BUF_X1 U127 ( .A(n1920), .Z(n6663) );
  BUF_X1 U128 ( .A(n1918), .Z(n6666) );
  BUF_X1 U129 ( .A(n1916), .Z(n6669) );
  BUF_X1 U130 ( .A(n1914), .Z(n6672) );
  BUF_X1 U131 ( .A(n1912), .Z(n6675) );
  BUF_X1 U132 ( .A(n1910), .Z(n6678) );
  BUF_X1 U133 ( .A(n1908), .Z(n6681) );
  BUF_X1 U134 ( .A(n1906), .Z(n6684) );
  BUF_X1 U135 ( .A(n1904), .Z(n6687) );
  BUF_X1 U136 ( .A(n1940), .Z(n6630) );
  BUF_X1 U137 ( .A(n1938), .Z(n6632) );
  BUF_X1 U138 ( .A(n1936), .Z(n6635) );
  BUF_X1 U139 ( .A(n1934), .Z(n6638) );
  BUF_X1 U140 ( .A(n1932), .Z(n6641) );
  BUF_X1 U141 ( .A(n1930), .Z(n6644) );
  BUF_X1 U142 ( .A(n1928), .Z(n6647) );
  BUF_X1 U143 ( .A(n1926), .Z(n6650) );
  BUF_X1 U144 ( .A(n1924), .Z(n6653) );
  BUF_X1 U145 ( .A(n1922), .Z(n6656) );
  BUF_X1 U146 ( .A(n1921), .Z(n6659) );
  BUF_X1 U147 ( .A(n1920), .Z(n6662) );
  BUF_X1 U148 ( .A(n1918), .Z(n6665) );
  BUF_X1 U149 ( .A(n1916), .Z(n6668) );
  BUF_X1 U150 ( .A(n1914), .Z(n6671) );
  BUF_X1 U151 ( .A(n1912), .Z(n6674) );
  BUF_X1 U152 ( .A(n1910), .Z(n6677) );
  BUF_X1 U153 ( .A(n1908), .Z(n6680) );
  BUF_X1 U154 ( .A(n1906), .Z(n6683) );
  BUF_X1 U155 ( .A(n1904), .Z(n6686) );
  BUF_X1 U156 ( .A(n1940), .Z(n6631) );
  BUF_X1 U157 ( .A(n1902), .Z(n6691) );
  BUF_X1 U158 ( .A(n1900), .Z(n6694) );
  BUF_X1 U159 ( .A(n1898), .Z(n6697) );
  BUF_X1 U160 ( .A(n1896), .Z(n6700) );
  BUF_X1 U161 ( .A(n1894), .Z(n6703) );
  BUF_X1 U162 ( .A(n1892), .Z(n6706) );
  BUF_X1 U163 ( .A(n1890), .Z(n6709) );
  BUF_X1 U164 ( .A(n1888), .Z(n6712) );
  BUF_X1 U165 ( .A(n1886), .Z(n6715) );
  BUF_X1 U166 ( .A(n1884), .Z(n6718) );
  BUF_X1 U167 ( .A(n1882), .Z(n6721) );
  BUF_X1 U168 ( .A(n1879), .Z(n6733) );
  BUF_X1 U169 ( .A(n1924), .Z(n6655) );
  BUF_X1 U170 ( .A(n1922), .Z(n6658) );
  BUF_X1 U171 ( .A(n1921), .Z(n6661) );
  BUF_X1 U172 ( .A(n1920), .Z(n6664) );
  BUF_X1 U173 ( .A(n1918), .Z(n6667) );
  BUF_X1 U174 ( .A(n1916), .Z(n6670) );
  BUF_X1 U175 ( .A(n1914), .Z(n6673) );
  BUF_X1 U176 ( .A(n1912), .Z(n6676) );
  BUF_X1 U177 ( .A(n1910), .Z(n6679) );
  BUF_X1 U178 ( .A(n1908), .Z(n6682) );
  BUF_X1 U179 ( .A(n1906), .Z(n6685) );
  BUF_X1 U180 ( .A(n1904), .Z(n6688) );
  BUF_X1 U181 ( .A(n1938), .Z(n6634) );
  BUF_X1 U182 ( .A(n1936), .Z(n6637) );
  BUF_X1 U183 ( .A(n1934), .Z(n6640) );
  BUF_X1 U184 ( .A(n1932), .Z(n6643) );
  BUF_X1 U185 ( .A(n1930), .Z(n6646) );
  BUF_X1 U186 ( .A(n1928), .Z(n6649) );
  BUF_X1 U187 ( .A(n1926), .Z(n6652) );
  INV_X1 U188 ( .A(n2368), .ZN(n6276) );
  INV_X1 U189 ( .A(n2369), .ZN(n6284) );
  INV_X1 U190 ( .A(n2375), .ZN(n6244) );
  INV_X1 U191 ( .A(n2376), .ZN(n6252) );
  INV_X1 U192 ( .A(n2368), .ZN(n6277) );
  INV_X1 U193 ( .A(n2375), .ZN(n6245) );
  AND2_X1 U194 ( .A1(n5080), .A2(n5045), .ZN(n2412) );
  INV_X1 U195 ( .A(n2354), .ZN(n6328) );
  INV_X1 U196 ( .A(n2355), .ZN(n6336) );
  INV_X1 U197 ( .A(n2361), .ZN(n6308) );
  INV_X1 U198 ( .A(n2362), .ZN(n6316) );
  INV_X1 U199 ( .A(n2355), .ZN(n6337) );
  INV_X1 U200 ( .A(n2362), .ZN(n6317) );
  INV_X1 U201 ( .A(n2386), .ZN(n6212) );
  INV_X1 U202 ( .A(n2387), .ZN(n6220) );
  INV_X1 U203 ( .A(n2407), .ZN(n6116) );
  INV_X1 U204 ( .A(n2393), .ZN(n6180) );
  INV_X1 U205 ( .A(n2394), .ZN(n6188) );
  INV_X1 U206 ( .A(n2400), .ZN(n6148) );
  INV_X1 U207 ( .A(n2401), .ZN(n6156) );
  INV_X1 U208 ( .A(n2408), .ZN(n6124) );
  INV_X1 U209 ( .A(n2387), .ZN(n6221) );
  INV_X1 U210 ( .A(n2408), .ZN(n6125) );
  INV_X1 U211 ( .A(n2394), .ZN(n6189) );
  INV_X1 U212 ( .A(n2401), .ZN(n6157) );
  BUF_X1 U213 ( .A(n6376), .Z(n6369) );
  BUF_X1 U214 ( .A(n6376), .Z(n6370) );
  BUF_X1 U215 ( .A(n6376), .Z(n6371) );
  BUF_X1 U216 ( .A(n6376), .Z(n6372) );
  BUF_X1 U217 ( .A(n6376), .Z(n6373) );
  BUF_X1 U218 ( .A(n6376), .Z(n6374) );
  BUF_X1 U219 ( .A(n6394), .Z(n6387) );
  BUF_X1 U220 ( .A(n6394), .Z(n6388) );
  BUF_X1 U221 ( .A(n6394), .Z(n6389) );
  BUF_X1 U222 ( .A(n6394), .Z(n6390) );
  BUF_X1 U223 ( .A(n6394), .Z(n6391) );
  BUF_X1 U224 ( .A(n6394), .Z(n6392) );
  BUF_X1 U225 ( .A(n6412), .Z(n6405) );
  BUF_X1 U226 ( .A(n6412), .Z(n6406) );
  BUF_X1 U227 ( .A(n6412), .Z(n6407) );
  BUF_X1 U228 ( .A(n6412), .Z(n6408) );
  BUF_X1 U229 ( .A(n6412), .Z(n6409) );
  BUF_X1 U230 ( .A(n6412), .Z(n6410) );
  BUF_X1 U231 ( .A(n6430), .Z(n6423) );
  BUF_X1 U232 ( .A(n6430), .Z(n6424) );
  BUF_X1 U233 ( .A(n6430), .Z(n6425) );
  BUF_X1 U234 ( .A(n6430), .Z(n6426) );
  BUF_X1 U235 ( .A(n6430), .Z(n6427) );
  BUF_X1 U236 ( .A(n6430), .Z(n6428) );
  BUF_X1 U237 ( .A(n6448), .Z(n6441) );
  BUF_X1 U238 ( .A(n6448), .Z(n6442) );
  BUF_X1 U239 ( .A(n6448), .Z(n6443) );
  BUF_X1 U240 ( .A(n6448), .Z(n6444) );
  BUF_X1 U241 ( .A(n6448), .Z(n6445) );
  BUF_X1 U242 ( .A(n6448), .Z(n6446) );
  BUF_X1 U243 ( .A(n6466), .Z(n6459) );
  BUF_X1 U244 ( .A(n6466), .Z(n6460) );
  BUF_X1 U245 ( .A(n6466), .Z(n6461) );
  BUF_X1 U246 ( .A(n6466), .Z(n6462) );
  BUF_X1 U247 ( .A(n6466), .Z(n6463) );
  BUF_X1 U248 ( .A(n6466), .Z(n6464) );
  BUF_X1 U249 ( .A(n6484), .Z(n6477) );
  BUF_X1 U250 ( .A(n6484), .Z(n6478) );
  BUF_X1 U251 ( .A(n6484), .Z(n6479) );
  BUF_X1 U252 ( .A(n6484), .Z(n6480) );
  BUF_X1 U253 ( .A(n6484), .Z(n6481) );
  BUF_X1 U254 ( .A(n6484), .Z(n6482) );
  BUF_X1 U255 ( .A(n6502), .Z(n6495) );
  BUF_X1 U256 ( .A(n6502), .Z(n6496) );
  BUF_X1 U257 ( .A(n6502), .Z(n6497) );
  BUF_X1 U258 ( .A(n6502), .Z(n6498) );
  BUF_X1 U259 ( .A(n6502), .Z(n6499) );
  BUF_X1 U260 ( .A(n6502), .Z(n6500) );
  BUF_X1 U261 ( .A(n6520), .Z(n6513) );
  BUF_X1 U262 ( .A(n6520), .Z(n6514) );
  BUF_X1 U263 ( .A(n6520), .Z(n6515) );
  BUF_X1 U264 ( .A(n6520), .Z(n6516) );
  BUF_X1 U265 ( .A(n6520), .Z(n6517) );
  BUF_X1 U266 ( .A(n6520), .Z(n6518) );
  BUF_X1 U267 ( .A(n6538), .Z(n6531) );
  BUF_X1 U268 ( .A(n6538), .Z(n6532) );
  BUF_X1 U269 ( .A(n6538), .Z(n6533) );
  BUF_X1 U270 ( .A(n6538), .Z(n6534) );
  BUF_X1 U271 ( .A(n6538), .Z(n6535) );
  BUF_X1 U272 ( .A(n6538), .Z(n6536) );
  BUF_X1 U273 ( .A(n6556), .Z(n6549) );
  BUF_X1 U274 ( .A(n6556), .Z(n6550) );
  BUF_X1 U275 ( .A(n6556), .Z(n6551) );
  BUF_X1 U276 ( .A(n6556), .Z(n6552) );
  BUF_X1 U277 ( .A(n6556), .Z(n6553) );
  BUF_X1 U278 ( .A(n6556), .Z(n6554) );
  BUF_X1 U279 ( .A(n6574), .Z(n6567) );
  BUF_X1 U280 ( .A(n6574), .Z(n6568) );
  BUF_X1 U281 ( .A(n6574), .Z(n6569) );
  BUF_X1 U282 ( .A(n6574), .Z(n6570) );
  BUF_X1 U283 ( .A(n6574), .Z(n6571) );
  BUF_X1 U284 ( .A(n6574), .Z(n6572) );
  BUF_X1 U285 ( .A(n6592), .Z(n6585) );
  BUF_X1 U286 ( .A(n6592), .Z(n6586) );
  BUF_X1 U287 ( .A(n6592), .Z(n6587) );
  BUF_X1 U288 ( .A(n6592), .Z(n6588) );
  BUF_X1 U289 ( .A(n6592), .Z(n6589) );
  BUF_X1 U290 ( .A(n6592), .Z(n6590) );
  BUF_X1 U291 ( .A(n6610), .Z(n6603) );
  BUF_X1 U292 ( .A(n6610), .Z(n6604) );
  BUF_X1 U293 ( .A(n6610), .Z(n6605) );
  BUF_X1 U294 ( .A(n6610), .Z(n6606) );
  BUF_X1 U295 ( .A(n6610), .Z(n6607) );
  BUF_X1 U296 ( .A(n6610), .Z(n6608) );
  BUF_X1 U297 ( .A(n6628), .Z(n6621) );
  BUF_X1 U298 ( .A(n6628), .Z(n6622) );
  BUF_X1 U299 ( .A(n6628), .Z(n6623) );
  BUF_X1 U300 ( .A(n6628), .Z(n6624) );
  BUF_X1 U301 ( .A(n6628), .Z(n6625) );
  BUF_X1 U302 ( .A(n6628), .Z(n6626) );
  BUF_X1 U303 ( .A(n6367), .Z(n6360) );
  BUF_X1 U304 ( .A(n6367), .Z(n6361) );
  BUF_X1 U305 ( .A(n6367), .Z(n6362) );
  BUF_X1 U306 ( .A(n6367), .Z(n6363) );
  BUF_X1 U307 ( .A(n6367), .Z(n6364) );
  BUF_X1 U308 ( .A(n6367), .Z(n6365) );
  BUF_X1 U309 ( .A(n6385), .Z(n6378) );
  BUF_X1 U310 ( .A(n6385), .Z(n6379) );
  BUF_X1 U311 ( .A(n6385), .Z(n6380) );
  BUF_X1 U312 ( .A(n6385), .Z(n6381) );
  BUF_X1 U313 ( .A(n6385), .Z(n6382) );
  BUF_X1 U314 ( .A(n6385), .Z(n6383) );
  BUF_X1 U315 ( .A(n6403), .Z(n6396) );
  BUF_X1 U316 ( .A(n6403), .Z(n6397) );
  BUF_X1 U317 ( .A(n6403), .Z(n6398) );
  BUF_X1 U318 ( .A(n6403), .Z(n6399) );
  BUF_X1 U319 ( .A(n6403), .Z(n6400) );
  BUF_X1 U320 ( .A(n6403), .Z(n6401) );
  BUF_X1 U321 ( .A(n6421), .Z(n6414) );
  BUF_X1 U322 ( .A(n6421), .Z(n6415) );
  BUF_X1 U323 ( .A(n6421), .Z(n6416) );
  BUF_X1 U324 ( .A(n6421), .Z(n6417) );
  BUF_X1 U325 ( .A(n6421), .Z(n6418) );
  BUF_X1 U326 ( .A(n6421), .Z(n6419) );
  BUF_X1 U327 ( .A(n6439), .Z(n6432) );
  BUF_X1 U328 ( .A(n6439), .Z(n6433) );
  BUF_X1 U329 ( .A(n6439), .Z(n6434) );
  BUF_X1 U330 ( .A(n6439), .Z(n6435) );
  BUF_X1 U331 ( .A(n6439), .Z(n6436) );
  BUF_X1 U332 ( .A(n6439), .Z(n6437) );
  BUF_X1 U333 ( .A(n6457), .Z(n6450) );
  BUF_X1 U334 ( .A(n6457), .Z(n6451) );
  BUF_X1 U335 ( .A(n6457), .Z(n6452) );
  BUF_X1 U336 ( .A(n6457), .Z(n6453) );
  BUF_X1 U337 ( .A(n6457), .Z(n6454) );
  BUF_X1 U338 ( .A(n6457), .Z(n6455) );
  BUF_X1 U339 ( .A(n6475), .Z(n6468) );
  BUF_X1 U340 ( .A(n6475), .Z(n6469) );
  BUF_X1 U341 ( .A(n6475), .Z(n6470) );
  BUF_X1 U342 ( .A(n6475), .Z(n6471) );
  BUF_X1 U343 ( .A(n6475), .Z(n6472) );
  BUF_X1 U344 ( .A(n6475), .Z(n6473) );
  BUF_X1 U345 ( .A(n6511), .Z(n6504) );
  BUF_X1 U346 ( .A(n6511), .Z(n6505) );
  BUF_X1 U347 ( .A(n6511), .Z(n6506) );
  BUF_X1 U348 ( .A(n6511), .Z(n6507) );
  BUF_X1 U349 ( .A(n6511), .Z(n6508) );
  BUF_X1 U350 ( .A(n6511), .Z(n6509) );
  BUF_X1 U351 ( .A(n6529), .Z(n6522) );
  BUF_X1 U352 ( .A(n6529), .Z(n6523) );
  BUF_X1 U353 ( .A(n6529), .Z(n6524) );
  BUF_X1 U354 ( .A(n6529), .Z(n6525) );
  BUF_X1 U355 ( .A(n6529), .Z(n6526) );
  BUF_X1 U356 ( .A(n6529), .Z(n6527) );
  BUF_X1 U357 ( .A(n6547), .Z(n6540) );
  BUF_X1 U358 ( .A(n6547), .Z(n6541) );
  BUF_X1 U359 ( .A(n6547), .Z(n6542) );
  BUF_X1 U360 ( .A(n6547), .Z(n6543) );
  BUF_X1 U361 ( .A(n6547), .Z(n6544) );
  BUF_X1 U362 ( .A(n6547), .Z(n6545) );
  BUF_X1 U363 ( .A(n6565), .Z(n6558) );
  BUF_X1 U364 ( .A(n6565), .Z(n6559) );
  BUF_X1 U365 ( .A(n6565), .Z(n6560) );
  BUF_X1 U366 ( .A(n6565), .Z(n6561) );
  BUF_X1 U367 ( .A(n6565), .Z(n6562) );
  BUF_X1 U368 ( .A(n6565), .Z(n6563) );
  BUF_X1 U369 ( .A(n6583), .Z(n6576) );
  BUF_X1 U370 ( .A(n6583), .Z(n6577) );
  BUF_X1 U371 ( .A(n6583), .Z(n6578) );
  BUF_X1 U372 ( .A(n6583), .Z(n6579) );
  BUF_X1 U373 ( .A(n6583), .Z(n6580) );
  BUF_X1 U374 ( .A(n6583), .Z(n6581) );
  BUF_X1 U375 ( .A(n6601), .Z(n6594) );
  BUF_X1 U376 ( .A(n6601), .Z(n6595) );
  BUF_X1 U377 ( .A(n6601), .Z(n6596) );
  BUF_X1 U378 ( .A(n6601), .Z(n6597) );
  BUF_X1 U379 ( .A(n6601), .Z(n6598) );
  BUF_X1 U380 ( .A(n6601), .Z(n6599) );
  BUF_X1 U381 ( .A(n6619), .Z(n6612) );
  BUF_X1 U382 ( .A(n6619), .Z(n6613) );
  BUF_X1 U383 ( .A(n6619), .Z(n6614) );
  BUF_X1 U384 ( .A(n6619), .Z(n6615) );
  BUF_X1 U385 ( .A(n6619), .Z(n6616) );
  BUF_X1 U386 ( .A(n6619), .Z(n6617) );
  BUF_X1 U387 ( .A(n6610), .Z(n6609) );
  BUF_X1 U388 ( .A(n6628), .Z(n6627) );
  BUF_X1 U389 ( .A(n6376), .Z(n6375) );
  BUF_X1 U390 ( .A(n6394), .Z(n6393) );
  BUF_X1 U391 ( .A(n6412), .Z(n6411) );
  BUF_X1 U392 ( .A(n6430), .Z(n6429) );
  BUF_X1 U393 ( .A(n6448), .Z(n6447) );
  BUF_X1 U394 ( .A(n6466), .Z(n6465) );
  BUF_X1 U395 ( .A(n6484), .Z(n6483) );
  BUF_X1 U396 ( .A(n6502), .Z(n6501) );
  BUF_X1 U397 ( .A(n6520), .Z(n6519) );
  BUF_X1 U398 ( .A(n6538), .Z(n6537) );
  BUF_X1 U399 ( .A(n6556), .Z(n6555) );
  BUF_X1 U400 ( .A(n6574), .Z(n6573) );
  BUF_X1 U401 ( .A(n6592), .Z(n6591) );
  BUF_X1 U402 ( .A(n6367), .Z(n6366) );
  BUF_X1 U403 ( .A(n6385), .Z(n6384) );
  BUF_X1 U404 ( .A(n6403), .Z(n6402) );
  BUF_X1 U405 ( .A(n6421), .Z(n6420) );
  BUF_X1 U406 ( .A(n6439), .Z(n6438) );
  BUF_X1 U407 ( .A(n6457), .Z(n6456) );
  BUF_X1 U408 ( .A(n6475), .Z(n6474) );
  BUF_X1 U409 ( .A(n6511), .Z(n6510) );
  BUF_X1 U410 ( .A(n6529), .Z(n6528) );
  BUF_X1 U411 ( .A(n6547), .Z(n6546) );
  BUF_X1 U412 ( .A(n6565), .Z(n6564) );
  BUF_X1 U413 ( .A(n6583), .Z(n6582) );
  BUF_X1 U414 ( .A(n6601), .Z(n6600) );
  BUF_X1 U415 ( .A(n6619), .Z(n6618) );
  INV_X1 U416 ( .A(n2160), .ZN(n6493) );
  OAI21_X1 U417 ( .B1(n1942), .B2(n2183), .A(RESET), .ZN(n2160) );
  INV_X1 U418 ( .A(n2346), .ZN(n6358) );
  NAND2_X1 U419 ( .A1(n5035), .A2(n5036), .ZN(OUT2[0]) );
  NOR4_X1 U420 ( .A1(n5063), .A2(n5064), .A3(n5065), .A4(n5066), .ZN(n5035) );
  NOR4_X1 U421 ( .A1(n5037), .A2(n5038), .A3(n5039), .A4(n5040), .ZN(n5036) );
  NAND2_X1 U422 ( .A1(n4661), .A2(n4662), .ZN(OUT2[1]) );
  NOR4_X1 U423 ( .A1(n4679), .A2(n4680), .A3(n4681), .A4(n4682), .ZN(n4661) );
  NOR4_X1 U424 ( .A1(n4663), .A2(n4664), .A3(n4665), .A4(n4666), .ZN(n4662) );
  NAND2_X1 U425 ( .A1(n3711), .A2(n3712), .ZN(OUT2[2]) );
  NOR4_X1 U426 ( .A1(n4305), .A2(n4306), .A3(n4307), .A4(n4308), .ZN(n3711) );
  NOR4_X1 U427 ( .A1(n3713), .A2(n3714), .A3(n3715), .A4(n3716), .ZN(n3712) );
  NAND2_X1 U428 ( .A1(n5001), .A2(n5002), .ZN(OUT2[10]) );
  NOR4_X1 U429 ( .A1(n5019), .A2(n5020), .A3(n5021), .A4(n5022), .ZN(n5001) );
  NOR4_X1 U430 ( .A1(n5003), .A2(n5004), .A3(n5005), .A4(n5006), .ZN(n5002) );
  NAND2_X1 U431 ( .A1(n4967), .A2(n4968), .ZN(OUT2[11]) );
  NOR4_X1 U432 ( .A1(n4985), .A2(n4986), .A3(n4987), .A4(n4988), .ZN(n4967) );
  NOR4_X1 U433 ( .A1(n4969), .A2(n4970), .A3(n4971), .A4(n4972), .ZN(n4968) );
  NAND2_X1 U434 ( .A1(n4933), .A2(n4934), .ZN(OUT2[12]) );
  NOR4_X1 U435 ( .A1(n4951), .A2(n4952), .A3(n4953), .A4(n4954), .ZN(n4933) );
  NOR4_X1 U436 ( .A1(n4935), .A2(n4936), .A3(n4937), .A4(n4938), .ZN(n4934) );
  NAND2_X1 U437 ( .A1(n4899), .A2(n4900), .ZN(OUT2[13]) );
  NOR4_X1 U438 ( .A1(n4917), .A2(n4918), .A3(n4919), .A4(n4920), .ZN(n4899) );
  NOR4_X1 U439 ( .A1(n4901), .A2(n4902), .A3(n4903), .A4(n4904), .ZN(n4900) );
  NAND2_X1 U440 ( .A1(n4865), .A2(n4866), .ZN(OUT2[14]) );
  NOR4_X1 U441 ( .A1(n4883), .A2(n4884), .A3(n4885), .A4(n4886), .ZN(n4865) );
  NOR4_X1 U442 ( .A1(n4867), .A2(n4868), .A3(n4869), .A4(n4870), .ZN(n4866) );
  NAND2_X1 U443 ( .A1(n4831), .A2(n4832), .ZN(OUT2[15]) );
  NOR4_X1 U444 ( .A1(n4849), .A2(n4850), .A3(n4851), .A4(n4852), .ZN(n4831) );
  NOR4_X1 U445 ( .A1(n4833), .A2(n4834), .A3(n4835), .A4(n4836), .ZN(n4832) );
  NAND2_X1 U446 ( .A1(n4797), .A2(n4798), .ZN(OUT2[16]) );
  NOR4_X1 U447 ( .A1(n4815), .A2(n4816), .A3(n4817), .A4(n4818), .ZN(n4797) );
  NOR4_X1 U448 ( .A1(n4799), .A2(n4800), .A3(n4801), .A4(n4802), .ZN(n4798) );
  NAND2_X1 U449 ( .A1(n4763), .A2(n4764), .ZN(OUT2[17]) );
  NOR4_X1 U450 ( .A1(n4781), .A2(n4782), .A3(n4783), .A4(n4784), .ZN(n4763) );
  NOR4_X1 U451 ( .A1(n4765), .A2(n4766), .A3(n4767), .A4(n4768), .ZN(n4764) );
  NAND2_X1 U452 ( .A1(n4729), .A2(n4730), .ZN(OUT2[18]) );
  NOR4_X1 U453 ( .A1(n4747), .A2(n4748), .A3(n4749), .A4(n4750), .ZN(n4729) );
  NOR4_X1 U454 ( .A1(n4731), .A2(n4732), .A3(n4733), .A4(n4734), .ZN(n4730) );
  NAND2_X1 U455 ( .A1(n4695), .A2(n4696), .ZN(OUT2[19]) );
  NOR4_X1 U456 ( .A1(n4713), .A2(n4714), .A3(n4715), .A4(n4716), .ZN(n4695) );
  NOR4_X1 U457 ( .A1(n4697), .A2(n4698), .A3(n4699), .A4(n4700), .ZN(n4696) );
  NAND2_X1 U458 ( .A1(n4627), .A2(n4628), .ZN(OUT2[20]) );
  NOR4_X1 U459 ( .A1(n4645), .A2(n4646), .A3(n4647), .A4(n4648), .ZN(n4627) );
  NOR4_X1 U460 ( .A1(n4629), .A2(n4630), .A3(n4631), .A4(n4632), .ZN(n4628) );
  NAND2_X1 U461 ( .A1(n4593), .A2(n4594), .ZN(OUT2[21]) );
  NOR4_X1 U462 ( .A1(n4611), .A2(n4612), .A3(n4613), .A4(n4614), .ZN(n4593) );
  NOR4_X1 U463 ( .A1(n4595), .A2(n4596), .A3(n4597), .A4(n4598), .ZN(n4594) );
  NAND2_X1 U464 ( .A1(n4559), .A2(n4560), .ZN(OUT2[22]) );
  NOR4_X1 U465 ( .A1(n4577), .A2(n4578), .A3(n4579), .A4(n4580), .ZN(n4559) );
  NOR4_X1 U466 ( .A1(n4561), .A2(n4562), .A3(n4563), .A4(n4564), .ZN(n4560) );
  NAND2_X1 U467 ( .A1(n4525), .A2(n4526), .ZN(OUT2[23]) );
  NOR4_X1 U468 ( .A1(n4543), .A2(n4544), .A3(n4545), .A4(n4546), .ZN(n4525) );
  NOR4_X1 U469 ( .A1(n4527), .A2(n4528), .A3(n4529), .A4(n4530), .ZN(n4526) );
  NAND2_X1 U470 ( .A1(n4491), .A2(n4492), .ZN(OUT2[24]) );
  NOR4_X1 U471 ( .A1(n4509), .A2(n4510), .A3(n4511), .A4(n4512), .ZN(n4491) );
  NOR4_X1 U472 ( .A1(n4493), .A2(n4494), .A3(n4495), .A4(n4496), .ZN(n4492) );
  NAND2_X1 U473 ( .A1(n4457), .A2(n4458), .ZN(OUT2[25]) );
  NOR4_X1 U474 ( .A1(n4475), .A2(n4476), .A3(n4477), .A4(n4478), .ZN(n4457) );
  NOR4_X1 U475 ( .A1(n4459), .A2(n4460), .A3(n4461), .A4(n4462), .ZN(n4458) );
  NAND2_X1 U476 ( .A1(n4423), .A2(n4424), .ZN(OUT2[26]) );
  NOR4_X1 U477 ( .A1(n4441), .A2(n4442), .A3(n4443), .A4(n4444), .ZN(n4423) );
  NOR4_X1 U478 ( .A1(n4425), .A2(n4426), .A3(n4427), .A4(n4428), .ZN(n4424) );
  NAND2_X1 U479 ( .A1(n4389), .A2(n4390), .ZN(OUT2[27]) );
  NOR4_X1 U480 ( .A1(n4407), .A2(n4408), .A3(n4409), .A4(n4410), .ZN(n4389) );
  NOR4_X1 U481 ( .A1(n4391), .A2(n4392), .A3(n4393), .A4(n4394), .ZN(n4390) );
  NAND2_X1 U482 ( .A1(n4355), .A2(n4356), .ZN(OUT2[28]) );
  NOR4_X1 U483 ( .A1(n4373), .A2(n4374), .A3(n4375), .A4(n4376), .ZN(n4355) );
  NOR4_X1 U484 ( .A1(n4357), .A2(n4358), .A3(n4359), .A4(n4360), .ZN(n4356) );
  NAND2_X1 U485 ( .A1(n4321), .A2(n4322), .ZN(OUT2[29]) );
  NOR4_X1 U486 ( .A1(n4339), .A2(n4340), .A3(n4341), .A4(n4342), .ZN(n4321) );
  NOR4_X1 U487 ( .A1(n4323), .A2(n4324), .A3(n4325), .A4(n4326), .ZN(n4322) );
  NAND2_X1 U488 ( .A1(n2652), .A2(n2653), .ZN(OUT2[30]) );
  NOR4_X1 U489 ( .A1(n3695), .A2(n3696), .A3(n3697), .A4(n3698), .ZN(n2652) );
  NOR4_X1 U490 ( .A1(n2654), .A2(n2655), .A3(n2656), .A4(n3682), .ZN(n2653) );
  NAND2_X1 U491 ( .A1(n2348), .A2(n2349), .ZN(OUT2[9]) );
  NOR4_X1 U492 ( .A1(n2382), .A2(n2383), .A3(n2384), .A4(n2385), .ZN(n2348) );
  NOR4_X1 U493 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(n2349) );
  NAND2_X1 U494 ( .A1(n2584), .A2(n2585), .ZN(OUT2[3]) );
  NOR4_X1 U495 ( .A1(n2602), .A2(n2603), .A3(n2604), .A4(n2605), .ZN(n2584) );
  NOR4_X1 U496 ( .A1(n2586), .A2(n2587), .A3(n2588), .A4(n2589), .ZN(n2585) );
  NAND2_X1 U497 ( .A1(n2550), .A2(n2551), .ZN(OUT2[4]) );
  NOR4_X1 U498 ( .A1(n2568), .A2(n2569), .A3(n2570), .A4(n2571), .ZN(n2550) );
  NOR4_X1 U499 ( .A1(n2552), .A2(n2553), .A3(n2554), .A4(n2555), .ZN(n2551) );
  NAND2_X1 U500 ( .A1(n2516), .A2(n2517), .ZN(OUT2[5]) );
  NOR4_X1 U501 ( .A1(n2534), .A2(n2535), .A3(n2536), .A4(n2537), .ZN(n2516) );
  NOR4_X1 U502 ( .A1(n2518), .A2(n2519), .A3(n2520), .A4(n2521), .ZN(n2517) );
  NAND2_X1 U503 ( .A1(n2482), .A2(n2483), .ZN(OUT2[6]) );
  NOR4_X1 U504 ( .A1(n2500), .A2(n2501), .A3(n2502), .A4(n2503), .ZN(n2482) );
  NOR4_X1 U505 ( .A1(n2484), .A2(n2485), .A3(n2486), .A4(n2487), .ZN(n2483) );
  NAND2_X1 U506 ( .A1(n2448), .A2(n2449), .ZN(OUT2[7]) );
  NOR4_X1 U507 ( .A1(n2466), .A2(n2467), .A3(n2468), .A4(n2469), .ZN(n2448) );
  NOR4_X1 U508 ( .A1(n2450), .A2(n2451), .A3(n2452), .A4(n2453), .ZN(n2449) );
  NAND2_X1 U509 ( .A1(n2414), .A2(n2415), .ZN(OUT2[8]) );
  NOR4_X1 U510 ( .A1(n2432), .A2(n2433), .A3(n2434), .A4(n2435), .ZN(n2414) );
  NOR4_X1 U511 ( .A1(n2416), .A2(n2417), .A3(n2418), .A4(n2419), .ZN(n2415) );
  NAND2_X1 U512 ( .A1(n2618), .A2(n2619), .ZN(OUT2[31]) );
  NOR4_X1 U513 ( .A1(n2636), .A2(n2637), .A3(n2638), .A4(n2639), .ZN(n2618) );
  NOR4_X1 U514 ( .A1(n2620), .A2(n2621), .A3(n2622), .A4(n2623), .ZN(n2619) );
  NOR3_X1 U515 ( .A1(n5692), .A2(n5691), .A3(n5705), .ZN(n5708) );
  AND2_X1 U516 ( .A1(n5686), .A2(n5689), .ZN(n6092) );
  AND2_X1 U517 ( .A1(n5686), .A2(n5689), .ZN(n6093) );
  AND2_X1 U518 ( .A1(n5686), .A2(n5685), .ZN(n6112) );
  AND2_X1 U519 ( .A1(n5686), .A2(n5685), .ZN(n6113) );
  AND2_X1 U520 ( .A1(n5684), .A2(n5689), .ZN(n6094) );
  AND2_X1 U521 ( .A1(n5684), .A2(n5689), .ZN(n6095) );
  AND2_X1 U522 ( .A1(n5684), .A2(n5685), .ZN(n6114) );
  AND2_X1 U523 ( .A1(n5684), .A2(n5685), .ZN(n6115) );
  AND2_X1 U524 ( .A1(n5686), .A2(n5689), .ZN(n5101) );
  AND2_X1 U525 ( .A1(n5686), .A2(n5685), .ZN(n5096) );
  AND2_X1 U526 ( .A1(n5684), .A2(n5689), .ZN(n5102) );
  AND2_X1 U527 ( .A1(n5684), .A2(n5685), .ZN(n5097) );
  NAND2_X1 U528 ( .A1(n5687), .A2(n5695), .ZN(n5103) );
  NAND2_X1 U529 ( .A1(n5687), .A2(n5694), .ZN(n5104) );
  NAND2_X1 U530 ( .A1(n5690), .A2(n5695), .ZN(n5108) );
  NAND2_X1 U531 ( .A1(n5690), .A2(n5694), .ZN(n5109) );
  OAI221_X1 U532 ( .B1(n2257), .B2(n5983), .C1(n2226), .C2(n5991), .A(n5475), 
        .ZN(n5474) );
  AOI22_X1 U533 ( .A1(n6003), .A2(n4650), .B1(n6008), .B2(n4651), .ZN(n5475)
         );
  OAI221_X1 U534 ( .B1(n2112), .B2(n6099), .C1(n2137), .C2(n6107), .A(n5467), 
        .ZN(n5466) );
  AOI22_X1 U535 ( .A1(n6112), .A2(n4634), .B1(n6114), .B2(n4635), .ZN(n5467)
         );
  OAI221_X1 U536 ( .B1(n2256), .B2(n5985), .C1(n2225), .C2(n5993), .A(n5457), 
        .ZN(n5456) );
  AOI22_X1 U537 ( .A1(n6003), .A2(n4616), .B1(n6009), .B2(n4617), .ZN(n5457)
         );
  OAI221_X1 U538 ( .B1(n2111), .B2(n6100), .C1(n2136), .C2(n6111), .A(n5449), 
        .ZN(n5448) );
  AOI22_X1 U539 ( .A1(n6113), .A2(n4600), .B1(n6115), .B2(n4601), .ZN(n5449)
         );
  OAI221_X1 U540 ( .B1(n2255), .B2(n5985), .C1(n2224), .C2(n5990), .A(n5439), 
        .ZN(n5438) );
  AOI22_X1 U541 ( .A1(n6001), .A2(n4582), .B1(n6010), .B2(n4583), .ZN(n5439)
         );
  OAI221_X1 U542 ( .B1(n2110), .B2(n6100), .C1(n2135), .C2(n6108), .A(n5431), 
        .ZN(n5430) );
  AOI22_X1 U543 ( .A1(n5096), .A2(n4566), .B1(n5097), .B2(n4567), .ZN(n5431)
         );
  OAI221_X1 U544 ( .B1(n2254), .B2(n5984), .C1(n2223), .C2(n5992), .A(n5421), 
        .ZN(n5420) );
  AOI22_X1 U545 ( .A1(n6002), .A2(n4548), .B1(n6011), .B2(n4549), .ZN(n5421)
         );
  OAI221_X1 U546 ( .B1(n2109), .B2(n6101), .C1(n2134), .C2(n6109), .A(n5413), 
        .ZN(n5412) );
  AOI22_X1 U547 ( .A1(n6112), .A2(n4532), .B1(n6114), .B2(n4533), .ZN(n5413)
         );
  OAI221_X1 U548 ( .B1(n2260), .B2(n5985), .C1(n2229), .C2(n5992), .A(n5547), 
        .ZN(n5546) );
  AOI22_X1 U549 ( .A1(n5999), .A2(n4786), .B1(n6008), .B2(n4787), .ZN(n5547)
         );
  OAI221_X1 U550 ( .B1(n2115), .B2(n6100), .C1(n2140), .C2(n6108), .A(n5539), 
        .ZN(n5538) );
  AOI22_X1 U551 ( .A1(n5096), .A2(n4770), .B1(n5097), .B2(n4771), .ZN(n5539)
         );
  OAI221_X1 U552 ( .B1(n2259), .B2(n5985), .C1(n2228), .C2(n5993), .A(n5529), 
        .ZN(n5528) );
  AOI22_X1 U553 ( .A1(n6000), .A2(n4752), .B1(n6007), .B2(n4753), .ZN(n5529)
         );
  OAI221_X1 U554 ( .B1(n2114), .B2(n6101), .C1(n2139), .C2(n6108), .A(n5521), 
        .ZN(n5520) );
  AOI22_X1 U555 ( .A1(n6112), .A2(n4736), .B1(n6114), .B2(n4737), .ZN(n5521)
         );
  OAI221_X1 U556 ( .B1(n2258), .B2(n5986), .C1(n2227), .C2(n5994), .A(n5511), 
        .ZN(n5510) );
  AOI22_X1 U557 ( .A1(n6001), .A2(n4718), .B1(n6010), .B2(n4719), .ZN(n5511)
         );
  OAI221_X1 U558 ( .B1(n2113), .B2(n6101), .C1(n2138), .C2(n6109), .A(n5503), 
        .ZN(n5502) );
  AOI22_X1 U559 ( .A1(n6113), .A2(n4702), .B1(n6115), .B2(n4703), .ZN(n5503)
         );
  OAI221_X1 U560 ( .B1(n2273), .B2(n5987), .C1(n2241), .C2(n5994), .A(n5493), 
        .ZN(n5492) );
  AOI22_X1 U561 ( .A1(n6002), .A2(n4684), .B1(n6011), .B2(n4685), .ZN(n5493)
         );
  OAI221_X1 U562 ( .B1(n2128), .B2(n6098), .C1(n2152), .C2(n6109), .A(n5485), 
        .ZN(n5484) );
  AOI22_X1 U563 ( .A1(n5096), .A2(n4668), .B1(n5097), .B2(n4669), .ZN(n5485)
         );
  OAI221_X1 U564 ( .B1(n2264), .B2(n5982), .C1(n2233), .C2(n5991), .A(n5619), 
        .ZN(n5618) );
  AOI22_X1 U565 ( .A1(n5998), .A2(n4922), .B1(n6006), .B2(n4923), .ZN(n5619)
         );
  OAI221_X1 U566 ( .B1(n2119), .B2(n6099), .C1(n2144), .C2(n6106), .A(n5611), 
        .ZN(n5610) );
  AOI22_X1 U567 ( .A1(n6113), .A2(n4906), .B1(n6115), .B2(n4907), .ZN(n5611)
         );
  OAI221_X1 U568 ( .B1(n2263), .B2(n5982), .C1(n2232), .C2(n5992), .A(n5601), 
        .ZN(n5600) );
  AOI22_X1 U569 ( .A1(n5998), .A2(n4888), .B1(n6007), .B2(n4889), .ZN(n5601)
         );
  OAI221_X1 U570 ( .B1(n2118), .B2(n6100), .C1(n2143), .C2(n6106), .A(n5593), 
        .ZN(n5592) );
  AOI22_X1 U571 ( .A1(n5096), .A2(n4872), .B1(n5097), .B2(n4873), .ZN(n5593)
         );
  OAI221_X1 U572 ( .B1(n2262), .B2(n5984), .C1(n2231), .C2(n5994), .A(n5583), 
        .ZN(n5582) );
  AOI22_X1 U573 ( .A1(n5999), .A2(n4854), .B1(n6008), .B2(n4855), .ZN(n5583)
         );
  OAI221_X1 U574 ( .B1(n2117), .B2(n6100), .C1(n2142), .C2(n6108), .A(n5575), 
        .ZN(n5574) );
  AOI22_X1 U575 ( .A1(n6112), .A2(n4838), .B1(n6114), .B2(n4839), .ZN(n5575)
         );
  OAI221_X1 U576 ( .B1(n2261), .B2(n5984), .C1(n2230), .C2(n5993), .A(n5565), 
        .ZN(n5564) );
  AOI22_X1 U577 ( .A1(n6003), .A2(n4820), .B1(n6009), .B2(n4821), .ZN(n5565)
         );
  OAI221_X1 U578 ( .B1(n2116), .B2(n6101), .C1(n2141), .C2(n6109), .A(n5557), 
        .ZN(n5556) );
  AOI22_X1 U579 ( .A1(n6113), .A2(n4804), .B1(n6115), .B2(n4805), .ZN(n5557)
         );
  OAI221_X1 U580 ( .B1(n2268), .B2(n5982), .C1(n2239), .C2(n5990), .A(n5187), 
        .ZN(n5186) );
  AOI22_X1 U581 ( .A1(n5999), .A2(n2505), .B1(n6008), .B2(n2506), .ZN(n5187)
         );
  OAI221_X1 U582 ( .B1(n2123), .B2(n6099), .C1(n2150), .C2(n6106), .A(n5179), 
        .ZN(n5178) );
  AOI22_X1 U583 ( .A1(n6113), .A2(n2489), .B1(n6115), .B2(n2490), .ZN(n5179)
         );
  OAI221_X1 U584 ( .B1(n2267), .B2(n5983), .C1(n2238), .C2(n5990), .A(n5169), 
        .ZN(n5168) );
  AOI22_X1 U585 ( .A1(n5999), .A2(n2471), .B1(n6009), .B2(n2472), .ZN(n5169)
         );
  OAI221_X1 U586 ( .B1(n2122), .B2(n6097), .C1(n2149), .C2(n6107), .A(n5161), 
        .ZN(n5160) );
  AOI22_X1 U587 ( .A1(n5096), .A2(n2455), .B1(n5097), .B2(n2456), .ZN(n5161)
         );
  OAI221_X1 U588 ( .B1(n2266), .B2(n5984), .C1(n2237), .C2(n5993), .A(n5151), 
        .ZN(n5150) );
  AOI22_X1 U589 ( .A1(n5999), .A2(n2437), .B1(n6009), .B2(n2438), .ZN(n5151)
         );
  OAI221_X1 U590 ( .B1(n2121), .B2(n6101), .C1(n2148), .C2(n6107), .A(n5143), 
        .ZN(n5142) );
  AOI22_X1 U591 ( .A1(n6112), .A2(n2421), .B1(n6114), .B2(n2422), .ZN(n5143)
         );
  OAI221_X1 U592 ( .B1(n2269), .B2(n5987), .C1(n2240), .C2(n5995), .A(n5205), 
        .ZN(n5204) );
  AOI22_X1 U593 ( .A1(n6002), .A2(n2539), .B1(n6007), .B2(n2540), .ZN(n5205)
         );
  OAI221_X1 U594 ( .B1(n2124), .B2(n6098), .C1(n2151), .C2(n6111), .A(n5197), 
        .ZN(n5196) );
  AOI22_X1 U595 ( .A1(n6112), .A2(n2523), .B1(n6114), .B2(n2524), .ZN(n5197)
         );
  OAI221_X1 U596 ( .B1(n2253), .B2(n5984), .C1(n2222), .C2(n5992), .A(n5403), 
        .ZN(n5402) );
  AOI22_X1 U597 ( .A1(n6003), .A2(n4514), .B1(n6010), .B2(n4515), .ZN(n5403)
         );
  OAI221_X1 U598 ( .B1(n2108), .B2(n6097), .C1(n2133), .C2(n6108), .A(n5395), 
        .ZN(n5394) );
  AOI22_X1 U599 ( .A1(n6113), .A2(n4498), .B1(n6115), .B2(n4499), .ZN(n5395)
         );
  OAI221_X1 U600 ( .B1(n2252), .B2(n5985), .C1(n2221), .C2(n5993), .A(n5385), 
        .ZN(n5384) );
  AOI22_X1 U601 ( .A1(n6003), .A2(n4480), .B1(n6009), .B2(n4481), .ZN(n5385)
         );
  OAI221_X1 U602 ( .B1(n2107), .B2(n6103), .C1(n2132), .C2(n6111), .A(n5377), 
        .ZN(n5376) );
  AOI22_X1 U603 ( .A1(n5096), .A2(n4464), .B1(n5097), .B2(n4465), .ZN(n5377)
         );
  OAI221_X1 U604 ( .B1(n2197), .B2(n5951), .C1(n2166), .C2(n5959), .A(n5476), 
        .ZN(n5473) );
  AOI22_X1 U605 ( .A1(n5971), .A2(n4653), .B1(n5976), .B2(n4654), .ZN(n5476)
         );
  OAI221_X1 U606 ( .B1(n2196), .B2(n5952), .C1(n2165), .C2(n5961), .A(n5458), 
        .ZN(n5455) );
  AOI22_X1 U607 ( .A1(n5971), .A2(n4619), .B1(n5977), .B2(n4620), .ZN(n5458)
         );
  OAI221_X1 U608 ( .B1(n2195), .B2(n5953), .C1(n2164), .C2(n5958), .A(n5440), 
        .ZN(n5437) );
  AOI22_X1 U609 ( .A1(n5969), .A2(n4585), .B1(n5978), .B2(n4586), .ZN(n5440)
         );
  OAI221_X1 U610 ( .B1(n2194), .B2(n5952), .C1(n2163), .C2(n5960), .A(n5422), 
        .ZN(n5419) );
  AOI22_X1 U611 ( .A1(n5970), .A2(n4551), .B1(n5979), .B2(n4552), .ZN(n5422)
         );
  OAI221_X1 U612 ( .B1(n2048), .B2(n6078), .C1(n2073), .C2(n6086), .A(n5414), 
        .ZN(n5411) );
  AOI22_X1 U613 ( .A1(n6092), .A2(n4535), .B1(n6094), .B2(n4536), .ZN(n5414)
         );
  OAI221_X1 U614 ( .B1(n2200), .B2(n5953), .C1(n2169), .C2(n5960), .A(n5548), 
        .ZN(n5545) );
  AOI22_X1 U615 ( .A1(n5967), .A2(n4789), .B1(n5976), .B2(n4790), .ZN(n5548)
         );
  OAI221_X1 U616 ( .B1(n2199), .B2(n5953), .C1(n2168), .C2(n5961), .A(n5530), 
        .ZN(n5527) );
  AOI22_X1 U617 ( .A1(n5968), .A2(n4755), .B1(n5975), .B2(n4756), .ZN(n5530)
         );
  OAI221_X1 U618 ( .B1(n2198), .B2(n5954), .C1(n2167), .C2(n5962), .A(n5512), 
        .ZN(n5509) );
  AOI22_X1 U619 ( .A1(n5969), .A2(n4721), .B1(n5978), .B2(n4722), .ZN(n5512)
         );
  OAI221_X1 U620 ( .B1(n2213), .B2(n5955), .C1(n2181), .C2(n5962), .A(n5494), 
        .ZN(n5491) );
  AOI22_X1 U621 ( .A1(n5970), .A2(n4687), .B1(n5979), .B2(n4688), .ZN(n5494)
         );
  OAI221_X1 U622 ( .B1(n2204), .B2(n5950), .C1(n2173), .C2(n5959), .A(n5620), 
        .ZN(n5617) );
  AOI22_X1 U623 ( .A1(n5966), .A2(n4925), .B1(n5974), .B2(n4926), .ZN(n5620)
         );
  OAI221_X1 U624 ( .B1(n2203), .B2(n5950), .C1(n2172), .C2(n5960), .A(n5602), 
        .ZN(n5599) );
  AOI22_X1 U625 ( .A1(n5966), .A2(n4891), .B1(n5975), .B2(n4892), .ZN(n5602)
         );
  OAI221_X1 U626 ( .B1(n2202), .B2(n5952), .C1(n2171), .C2(n5962), .A(n5584), 
        .ZN(n5581) );
  AOI22_X1 U627 ( .A1(n5967), .A2(n4857), .B1(n5976), .B2(n4858), .ZN(n5584)
         );
  OAI221_X1 U628 ( .B1(n2201), .B2(n5952), .C1(n2170), .C2(n5961), .A(n5566), 
        .ZN(n5563) );
  AOI22_X1 U629 ( .A1(n5971), .A2(n4823), .B1(n5977), .B2(n4824), .ZN(n5566)
         );
  OAI221_X1 U630 ( .B1(n2208), .B2(n5950), .C1(n2179), .C2(n5958), .A(n5188), 
        .ZN(n5185) );
  AOI22_X1 U631 ( .A1(n5967), .A2(n2508), .B1(n5976), .B2(n2509), .ZN(n5188)
         );
  OAI221_X1 U632 ( .B1(n2207), .B2(n5951), .C1(n2178), .C2(n5958), .A(n5170), 
        .ZN(n5167) );
  AOI22_X1 U633 ( .A1(n5967), .A2(n2474), .B1(n5977), .B2(n2475), .ZN(n5170)
         );
  OAI221_X1 U634 ( .B1(n2206), .B2(n5952), .C1(n2177), .C2(n5961), .A(n5152), 
        .ZN(n5149) );
  AOI22_X1 U635 ( .A1(n5967), .A2(n2440), .B1(n5977), .B2(n2441), .ZN(n5152)
         );
  OAI221_X1 U636 ( .B1(n2059), .B2(n6079), .C1(n2087), .C2(n6087), .A(n5100), 
        .ZN(n5091) );
  AOI22_X1 U637 ( .A1(n6093), .A2(n2365), .B1(n6095), .B2(n2367), .ZN(n5100)
         );
  OAI221_X1 U638 ( .B1(n2209), .B2(n5955), .C1(n2180), .C2(n5963), .A(n5206), 
        .ZN(n5203) );
  AOI22_X1 U639 ( .A1(n5970), .A2(n2542), .B1(n5975), .B2(n2543), .ZN(n5206)
         );
  OAI221_X1 U640 ( .B1(n2193), .B2(n5953), .C1(n2162), .C2(n5960), .A(n5404), 
        .ZN(n5401) );
  AOI22_X1 U641 ( .A1(n5971), .A2(n4517), .B1(n5978), .B2(n4518), .ZN(n5404)
         );
  OAI221_X1 U642 ( .B1(n2192), .B2(n5953), .C1(n2161), .C2(n5961), .A(n5386), 
        .ZN(n5383) );
  AOI22_X1 U643 ( .A1(n5971), .A2(n4483), .B1(n5977), .B2(n4484), .ZN(n5386)
         );
  OAI221_X1 U644 ( .B1(n2291), .B2(n5918), .C1(n2316), .C2(n5926), .A(n5477), 
        .ZN(n5472) );
  AOI22_X1 U645 ( .A1(n5939), .A2(n4656), .B1(n5944), .B2(n4657), .ZN(n5477)
         );
  OAI221_X1 U646 ( .B1(n1990), .B2(n6045), .C1(n2016), .C2(n6053), .A(n5469), 
        .ZN(n5464) );
  AOI22_X1 U647 ( .A1(n6067), .A2(n4640), .B1(n6074), .B2(n4641), .ZN(n5469)
         );
  OAI221_X1 U648 ( .B1(n2290), .B2(n5922), .C1(n2315), .C2(n5927), .A(n5459), 
        .ZN(n5454) );
  AOI22_X1 U649 ( .A1(n5939), .A2(n4622), .B1(n5945), .B2(n4623), .ZN(n5459)
         );
  OAI221_X1 U650 ( .B1(n1989), .B2(n6047), .C1(n2015), .C2(n6056), .A(n5451), 
        .ZN(n5446) );
  AOI22_X1 U651 ( .A1(n6067), .A2(n4606), .B1(n6074), .B2(n4607), .ZN(n5451)
         );
  OAI221_X1 U652 ( .B1(n2289), .B2(n5920), .C1(n2314), .C2(n5928), .A(n5441), 
        .ZN(n5436) );
  AOI22_X1 U653 ( .A1(n5937), .A2(n4588), .B1(n5946), .B2(n4589), .ZN(n5441)
         );
  OAI221_X1 U654 ( .B1(n1988), .B2(n6048), .C1(n2014), .C2(n6059), .A(n5433), 
        .ZN(n5428) );
  AOI22_X1 U655 ( .A1(n6065), .A2(n4572), .B1(n6073), .B2(n4573), .ZN(n5433)
         );
  OAI221_X1 U656 ( .B1(n2288), .B2(n5921), .C1(n2313), .C2(n5929), .A(n5423), 
        .ZN(n5418) );
  AOI22_X1 U657 ( .A1(n5938), .A2(n4554), .B1(n5947), .B2(n4555), .ZN(n5423)
         );
  OAI221_X1 U658 ( .B1(n1987), .B2(n6047), .C1(n2013), .C2(n6055), .A(n5415), 
        .ZN(n5410) );
  AOI22_X1 U659 ( .A1(n6066), .A2(n4538), .B1(n6073), .B2(n4539), .ZN(n5415)
         );
  OAI221_X1 U660 ( .B1(n2294), .B2(n5920), .C1(n2319), .C2(n5928), .A(n5549), 
        .ZN(n5544) );
  AOI22_X1 U661 ( .A1(n5935), .A2(n4792), .B1(n5944), .B2(n4793), .ZN(n5549)
         );
  OAI221_X1 U662 ( .B1(n1993), .B2(n6047), .C1(n2019), .C2(n6055), .A(n5541), 
        .ZN(n5536) );
  AOI22_X1 U663 ( .A1(n6063), .A2(n4776), .B1(n6074), .B2(n4777), .ZN(n5541)
         );
  OAI221_X1 U664 ( .B1(n2293), .B2(n5920), .C1(n2318), .C2(n5928), .A(n5531), 
        .ZN(n5526) );
  AOI22_X1 U665 ( .A1(n5936), .A2(n4758), .B1(n5943), .B2(n4759), .ZN(n5531)
         );
  OAI221_X1 U666 ( .B1(n1992), .B2(n6049), .C1(n2018), .C2(n6058), .A(n5523), 
        .ZN(n5518) );
  AOI22_X1 U667 ( .A1(n6064), .A2(n4742), .B1(n6075), .B2(n4743), .ZN(n5523)
         );
  OAI221_X1 U668 ( .B1(n2292), .B2(n5922), .C1(n2317), .C2(n5930), .A(n5513), 
        .ZN(n5508) );
  AOI22_X1 U669 ( .A1(n5937), .A2(n4724), .B1(n5946), .B2(n4725), .ZN(n5513)
         );
  OAI221_X1 U670 ( .B1(n1991), .B2(n6049), .C1(n2017), .C2(n6056), .A(n5505), 
        .ZN(n5500) );
  AOI22_X1 U671 ( .A1(n6065), .A2(n4708), .B1(n6073), .B2(n4709), .ZN(n5505)
         );
  OAI221_X1 U672 ( .B1(n2307), .B2(n5923), .C1(n2331), .C2(n5929), .A(n5495), 
        .ZN(n5490) );
  AOI22_X1 U673 ( .A1(n5938), .A2(n4690), .B1(n5947), .B2(n4691), .ZN(n5495)
         );
  OAI221_X1 U674 ( .B1(n2007), .B2(n6050), .C1(n2032), .C2(n6057), .A(n5487), 
        .ZN(n5482) );
  AOI22_X1 U675 ( .A1(n6066), .A2(n4674), .B1(n6073), .B2(n4675), .ZN(n5487)
         );
  OAI221_X1 U676 ( .B1(n2298), .B2(n5919), .C1(n2323), .C2(n5925), .A(n5621), 
        .ZN(n5616) );
  AOI22_X1 U677 ( .A1(n5934), .A2(n4928), .B1(n5942), .B2(n4929), .ZN(n5621)
         );
  OAI221_X1 U678 ( .B1(n1997), .B2(n6046), .C1(n2023), .C2(n6054), .A(n5613), 
        .ZN(n5608) );
  AOI22_X1 U679 ( .A1(n6062), .A2(n4912), .B1(n6071), .B2(n4913), .ZN(n5613)
         );
  OAI221_X1 U680 ( .B1(n2297), .B2(n5921), .C1(n2322), .C2(n5927), .A(n5603), 
        .ZN(n5598) );
  AOI22_X1 U681 ( .A1(n5934), .A2(n4894), .B1(n5943), .B2(n4895), .ZN(n5603)
         );
  OAI221_X1 U682 ( .B1(n1996), .B2(n6047), .C1(n2022), .C2(n6055), .A(n5595), 
        .ZN(n5590) );
  AOI22_X1 U683 ( .A1(n6062), .A2(n4878), .B1(n6071), .B2(n4879), .ZN(n5595)
         );
  OAI221_X1 U684 ( .B1(n2296), .B2(n5920), .C1(n2321), .C2(n5928), .A(n5585), 
        .ZN(n5580) );
  AOI22_X1 U685 ( .A1(n5935), .A2(n4860), .B1(n5944), .B2(n4861), .ZN(n5585)
         );
  OAI221_X1 U686 ( .B1(n1995), .B2(n6048), .C1(n2021), .C2(n6057), .A(n5577), 
        .ZN(n5572) );
  AOI22_X1 U687 ( .A1(n6063), .A2(n4844), .B1(n6072), .B2(n4845), .ZN(n5577)
         );
  OAI221_X1 U688 ( .B1(n2295), .B2(n5921), .C1(n2320), .C2(n5929), .A(n5567), 
        .ZN(n5562) );
  AOI22_X1 U689 ( .A1(n5939), .A2(n4826), .B1(n5945), .B2(n4827), .ZN(n5567)
         );
  OAI221_X1 U690 ( .B1(n1994), .B2(n6048), .C1(n2020), .C2(n6055), .A(n5559), 
        .ZN(n5554) );
  AOI22_X1 U691 ( .A1(n6067), .A2(n4810), .B1(n6072), .B2(n4811), .ZN(n5559)
         );
  OAI221_X1 U692 ( .B1(n1998), .B2(n6046), .C1(n2024), .C2(n6054), .A(n5631), 
        .ZN(n5626) );
  AOI22_X1 U693 ( .A1(n6066), .A2(n4946), .B1(n6072), .B2(n4947), .ZN(n5631)
         );
  OAI221_X1 U694 ( .B1(n2302), .B2(n5918), .C1(n2329), .C2(n5925), .A(n5189), 
        .ZN(n5184) );
  AOI22_X1 U695 ( .A1(n5935), .A2(n2511), .B1(n5944), .B2(n2512), .ZN(n5189)
         );
  OAI221_X1 U696 ( .B1(n2002), .B2(n6045), .C1(n2029), .C2(n6053), .A(n5181), 
        .ZN(n5176) );
  AOI22_X1 U697 ( .A1(n6063), .A2(n2495), .B1(n6072), .B2(n2496), .ZN(n5181)
         );
  OAI221_X1 U698 ( .B1(n2301), .B2(n5918), .C1(n2328), .C2(n5926), .A(n5171), 
        .ZN(n5166) );
  AOI22_X1 U699 ( .A1(n5935), .A2(n2477), .B1(n5945), .B2(n2478), .ZN(n5171)
         );
  OAI221_X1 U700 ( .B1(n2001), .B2(n6051), .C1(n2028), .C2(n6053), .A(n5163), 
        .ZN(n5158) );
  AOI22_X1 U701 ( .A1(n6063), .A2(n2461), .B1(n6072), .B2(n2462), .ZN(n5163)
         );
  OAI221_X1 U702 ( .B1(n2300), .B2(n5919), .C1(n2327), .C2(n5925), .A(n5153), 
        .ZN(n5148) );
  AOI22_X1 U703 ( .A1(n5935), .A2(n2443), .B1(n5945), .B2(n2444), .ZN(n5153)
         );
  OAI221_X1 U704 ( .B1(n1999), .B2(n6046), .C1(n2027), .C2(n6054), .A(n5105), 
        .ZN(n5090) );
  AOI22_X1 U705 ( .A1(n6064), .A2(n2372), .B1(n6073), .B2(n2374), .ZN(n5105)
         );
  OAI221_X1 U706 ( .B1(n2004), .B2(n6051), .C1(n2031), .C2(n6058), .A(n5217), 
        .ZN(n5212) );
  AOI22_X1 U707 ( .A1(n6066), .A2(n2563), .B1(n6071), .B2(n2564), .ZN(n5217)
         );
  OAI221_X1 U708 ( .B1(n2303), .B2(n5923), .C1(n2330), .C2(n5931), .A(n5207), 
        .ZN(n5202) );
  AOI22_X1 U709 ( .A1(n5938), .A2(n2545), .B1(n5943), .B2(n2546), .ZN(n5207)
         );
  OAI221_X1 U710 ( .B1(n2003), .B2(n6050), .C1(n2030), .C2(n6059), .A(n5199), 
        .ZN(n5194) );
  AOI22_X1 U711 ( .A1(n6062), .A2(n2529), .B1(n6071), .B2(n2530), .ZN(n5199)
         );
  OAI221_X1 U712 ( .B1(n2287), .B2(n5921), .C1(n2312), .C2(n5927), .A(n5405), 
        .ZN(n5400) );
  AOI22_X1 U713 ( .A1(n5939), .A2(n4520), .B1(n5946), .B2(n4521), .ZN(n5405)
         );
  OAI221_X1 U714 ( .B1(n1986), .B2(n6048), .C1(n2012), .C2(n6055), .A(n5397), 
        .ZN(n5392) );
  AOI22_X1 U715 ( .A1(n6067), .A2(n4504), .B1(n6074), .B2(n4505), .ZN(n5397)
         );
  OAI221_X1 U716 ( .B1(n2286), .B2(n5921), .C1(n2311), .C2(n5927), .A(n5387), 
        .ZN(n5382) );
  AOI22_X1 U717 ( .A1(n5939), .A2(n4486), .B1(n5945), .B2(n4487), .ZN(n5387)
         );
  OAI221_X1 U718 ( .B1(n1985), .B2(n6048), .C1(n2011), .C2(n6059), .A(n5379), 
        .ZN(n5374) );
  AOI22_X1 U719 ( .A1(n6067), .A2(n4470), .B1(n6075), .B2(n4471), .ZN(n5379)
         );
  OAI221_X1 U720 ( .B1(n1903), .B2(n6015), .C1(n1949), .C2(n6024), .A(n5470), 
        .ZN(n5463) );
  AOI22_X1 U721 ( .A1(n6035), .A2(n4643), .B1(n6040), .B2(n4644), .ZN(n5470)
         );
  OAI221_X1 U722 ( .B1(n1901), .B2(n6015), .C1(n1948), .C2(n6023), .A(n5452), 
        .ZN(n5445) );
  AOI22_X1 U723 ( .A1(n6035), .A2(n4609), .B1(n6041), .B2(n4610), .ZN(n5452)
         );
  OAI221_X1 U724 ( .B1(n1899), .B2(n6016), .C1(n1947), .C2(n6024), .A(n5434), 
        .ZN(n5427) );
  AOI22_X1 U725 ( .A1(n6033), .A2(n4575), .B1(n6042), .B2(n4576), .ZN(n5434)
         );
  OAI221_X1 U726 ( .B1(n1909), .B2(n6015), .C1(n1952), .C2(n6024), .A(n5542), 
        .ZN(n5535) );
  AOI22_X1 U727 ( .A1(n6032), .A2(n4779), .B1(n6040), .B2(n4780), .ZN(n5542)
         );
  OAI221_X1 U728 ( .B1(n1907), .B2(n6017), .C1(n1951), .C2(n6027), .A(n5524), 
        .ZN(n5517) );
  AOI22_X1 U729 ( .A1(n6034), .A2(n4745), .B1(n6039), .B2(n4746), .ZN(n5524)
         );
  OAI221_X1 U730 ( .B1(n1905), .B2(n6017), .C1(n1950), .C2(n6022), .A(n5506), 
        .ZN(n5499) );
  AOI22_X1 U731 ( .A1(n6033), .A2(n4711), .B1(n6042), .B2(n4712), .ZN(n5506)
         );
  OAI221_X1 U732 ( .B1(n1939), .B2(n6019), .C1(n1965), .C2(n6025), .A(n5488), 
        .ZN(n5481) );
  AOI22_X1 U733 ( .A1(n6034), .A2(n4677), .B1(n6043), .B2(n4678), .ZN(n5488)
         );
  OAI221_X1 U734 ( .B1(n1917), .B2(n6016), .C1(n1956), .C2(n6021), .A(n5614), 
        .ZN(n5607) );
  AOI22_X1 U735 ( .A1(n6031), .A2(n4915), .B1(n6038), .B2(n4916), .ZN(n5614)
         );
  OAI221_X1 U736 ( .B1(n1915), .B2(n6015), .C1(n1955), .C2(n6023), .A(n5596), 
        .ZN(n5589) );
  AOI22_X1 U737 ( .A1(n6031), .A2(n4881), .B1(n6039), .B2(n4882), .ZN(n5596)
         );
  OAI221_X1 U738 ( .B1(n1913), .B2(n6016), .C1(n1954), .C2(n6024), .A(n5578), 
        .ZN(n5571) );
  AOI22_X1 U739 ( .A1(n6032), .A2(n4847), .B1(n6040), .B2(n4848), .ZN(n5578)
         );
  OAI221_X1 U740 ( .B1(n1911), .B2(n6014), .C1(n1953), .C2(n6022), .A(n5560), 
        .ZN(n5553) );
  AOI22_X1 U741 ( .A1(n6033), .A2(n4813), .B1(n6041), .B2(n4814), .ZN(n5560)
         );
  OAI221_X1 U742 ( .B1(n1929), .B2(n6015), .C1(n1962), .C2(n6021), .A(n5182), 
        .ZN(n5175) );
  AOI22_X1 U743 ( .A1(n6032), .A2(n2498), .B1(n6040), .B2(n2499), .ZN(n5182)
         );
  OAI221_X1 U744 ( .B1(n1927), .B2(n6014), .C1(n1961), .C2(n6027), .A(n5164), 
        .ZN(n5157) );
  AOI22_X1 U745 ( .A1(n6031), .A2(n2464), .B1(n6041), .B2(n2465), .ZN(n5164)
         );
  OAI221_X1 U746 ( .B1(n1933), .B2(n6018), .C1(n1964), .C2(n6027), .A(n5218), 
        .ZN(n5211) );
  AOI22_X1 U747 ( .A1(n6033), .A2(n2566), .B1(n6038), .B2(n2567), .ZN(n5218)
         );
  OAI221_X1 U748 ( .B1(n1931), .B2(n6019), .C1(n1963), .C2(n6025), .A(n5200), 
        .ZN(n5193) );
  AOI22_X1 U749 ( .A1(n6031), .A2(n2532), .B1(n6039), .B2(n2533), .ZN(n5200)
         );
  OAI221_X1 U750 ( .B1(n1895), .B2(n6016), .C1(n1945), .C2(n6023), .A(n5398), 
        .ZN(n5391) );
  AOI22_X1 U751 ( .A1(n6035), .A2(n4507), .B1(n6042), .B2(n4508), .ZN(n5398)
         );
  NAND2_X1 U752 ( .A1(n5686), .A2(n5687), .ZN(n5093) );
  NAND2_X1 U753 ( .A1(n5684), .A2(n5687), .ZN(n5094) );
  NAND2_X1 U754 ( .A1(n5686), .A2(n5690), .ZN(n5098) );
  NAND2_X1 U755 ( .A1(n5684), .A2(n5690), .ZN(n5099) );
  NAND2_X1 U756 ( .A1(n5703), .A2(n5687), .ZN(n5117) );
  NAND2_X1 U757 ( .A1(n5702), .A2(n5687), .ZN(n5118) );
  NAND2_X1 U758 ( .A1(n5703), .A2(n5690), .ZN(n5122) );
  NAND2_X1 U759 ( .A1(n5702), .A2(n5690), .ZN(n5123) );
  NAND2_X1 U760 ( .A1(n5707), .A2(n5690), .ZN(n5127) );
  NAND2_X1 U761 ( .A1(n5708), .A2(n5690), .ZN(n5128) );
  NAND2_X1 U762 ( .A1(n5708), .A2(n5687), .ZN(n5132) );
  NAND2_X1 U763 ( .A1(n5707), .A2(n5687), .ZN(n5133) );
  AOI22_X1 U764 ( .A1(n6092), .A2(n4637), .B1(n6094), .B2(n4638), .ZN(n5468)
         );
  AOI22_X1 U765 ( .A1(n6093), .A2(n4603), .B1(n6095), .B2(n4604), .ZN(n5450)
         );
  AOI22_X1 U766 ( .A1(n5101), .A2(n4569), .B1(n5102), .B2(n4570), .ZN(n5432)
         );
  AOI22_X1 U767 ( .A1(n6034), .A2(n4541), .B1(n6043), .B2(n4542), .ZN(n5416)
         );
  AOI22_X1 U768 ( .A1(n5101), .A2(n4773), .B1(n5102), .B2(n4774), .ZN(n5540)
         );
  AOI22_X1 U769 ( .A1(n6092), .A2(n4739), .B1(n6094), .B2(n4740), .ZN(n5522)
         );
  AOI22_X1 U770 ( .A1(n6093), .A2(n4705), .B1(n6095), .B2(n4706), .ZN(n5504)
         );
  AOI22_X1 U771 ( .A1(n5101), .A2(n4671), .B1(n5102), .B2(n4672), .ZN(n5486)
         );
  AOI22_X1 U772 ( .A1(n6093), .A2(n4909), .B1(n6095), .B2(n4910), .ZN(n5612)
         );
  AOI22_X1 U773 ( .A1(n5101), .A2(n4875), .B1(n5102), .B2(n4876), .ZN(n5594)
         );
  AOI22_X1 U774 ( .A1(n6092), .A2(n4841), .B1(n6094), .B2(n4842), .ZN(n5576)
         );
  AOI22_X1 U775 ( .A1(n6093), .A2(n4807), .B1(n6095), .B2(n4808), .ZN(n5558)
         );
  AOI22_X1 U776 ( .A1(n6092), .A2(n5049), .B1(n6094), .B2(n5050), .ZN(n5688)
         );
  AOI22_X1 U777 ( .A1(n6093), .A2(n5011), .B1(n6095), .B2(n5012), .ZN(n5666)
         );
  AOI22_X1 U778 ( .A1(n5101), .A2(n4977), .B1(n5102), .B2(n4978), .ZN(n5648)
         );
  AOI22_X1 U779 ( .A1(n6034), .A2(n4949), .B1(n6038), .B2(n4950), .ZN(n5632)
         );
  AOI22_X1 U780 ( .A1(n6093), .A2(n2492), .B1(n6095), .B2(n2493), .ZN(n5180)
         );
  AOI22_X1 U781 ( .A1(n5101), .A2(n2458), .B1(n5102), .B2(n2459), .ZN(n5162)
         );
  AOI22_X1 U782 ( .A1(n6092), .A2(n2424), .B1(n6094), .B2(n2425), .ZN(n5144)
         );
  AOI22_X1 U783 ( .A1(n6032), .A2(n2379), .B1(n6042), .B2(n2381), .ZN(n5110)
         );
  AOI22_X1 U784 ( .A1(n6092), .A2(n2628), .B1(n6094), .B2(n2629), .ZN(n5252)
         );
  AOI22_X1 U785 ( .A1(n6093), .A2(n2594), .B1(n6095), .B2(n2595), .ZN(n5234)
         );
  AOI22_X1 U786 ( .A1(n5101), .A2(n2560), .B1(n5102), .B2(n2561), .ZN(n5216)
         );
  AOI22_X1 U787 ( .A1(n6092), .A2(n2526), .B1(n6094), .B2(n2527), .ZN(n5198)
         );
  AOI22_X1 U788 ( .A1(n6093), .A2(n4501), .B1(n6095), .B2(n4502), .ZN(n5396)
         );
  AOI22_X1 U789 ( .A1(n5101), .A2(n4467), .B1(n5102), .B2(n4468), .ZN(n5378)
         );
  AOI22_X1 U790 ( .A1(n6035), .A2(n4439), .B1(n6043), .B2(n4440), .ZN(n5362)
         );
  AOI22_X1 U791 ( .A1(n6034), .A2(n4405), .B1(n6043), .B2(n4406), .ZN(n5344)
         );
  AOI22_X1 U792 ( .A1(n6033), .A2(n4371), .B1(n6038), .B2(n4372), .ZN(n5326)
         );
  AOI22_X1 U793 ( .A1(n6033), .A2(n4337), .B1(n6039), .B2(n4338), .ZN(n5308)
         );
  AOI22_X1 U794 ( .A1(n6093), .A2(n3721), .B1(n6095), .B2(n4298), .ZN(n5288)
         );
  AOI22_X1 U795 ( .A1(n5101), .A2(n3687), .B1(n5102), .B2(n3688), .ZN(n5270)
         );
  AND2_X1 U796 ( .A1(n5689), .A2(n5695), .ZN(n5111) );
  AND2_X1 U797 ( .A1(n5685), .A2(n5694), .ZN(n5107) );
  AND2_X1 U798 ( .A1(n5685), .A2(n5695), .ZN(n5106) );
  AND2_X1 U799 ( .A1(n5702), .A2(n5689), .ZN(n5126) );
  AND2_X1 U800 ( .A1(n5703), .A2(n5689), .ZN(n5125) );
  AND2_X1 U801 ( .A1(n5707), .A2(n5689), .ZN(n5131) );
  AND2_X1 U802 ( .A1(n5708), .A2(n5689), .ZN(n5130) );
  AND2_X1 U803 ( .A1(n5694), .A2(n5689), .ZN(n5112) );
  AND2_X1 U804 ( .A1(n5702), .A2(n5685), .ZN(n5121) );
  AND2_X1 U805 ( .A1(n5703), .A2(n5685), .ZN(n5120) );
  AND2_X1 U806 ( .A1(n5707), .A2(n5685), .ZN(n5135) );
  NAND2_X1 U807 ( .A1(n5461), .A2(n5462), .ZN(OUT1[20]) );
  NOR4_X1 U808 ( .A1(n5463), .A2(n5464), .A3(n5465), .A4(n5466), .ZN(n5462) );
  NOR4_X1 U809 ( .A1(n5471), .A2(n5472), .A3(n5473), .A4(n5474), .ZN(n5461) );
  OAI221_X1 U810 ( .B1(n2051), .B2(n6083), .C1(n2076), .C2(n6088), .A(n5468), 
        .ZN(n5465) );
  NAND2_X1 U811 ( .A1(n5533), .A2(n5534), .ZN(OUT1[17]) );
  NOR4_X1 U812 ( .A1(n5535), .A2(n5536), .A3(n5537), .A4(n5538), .ZN(n5534) );
  NOR4_X1 U813 ( .A1(n5543), .A2(n5544), .A3(n5545), .A4(n5546), .ZN(n5533) );
  OAI221_X1 U814 ( .B1(n2054), .B2(n6081), .C1(n2079), .C2(n6088), .A(n5540), 
        .ZN(n5537) );
  NAND2_X1 U815 ( .A1(n5605), .A2(n5606), .ZN(OUT1[13]) );
  NOR4_X1 U816 ( .A1(n5607), .A2(n5608), .A3(n5609), .A4(n5610), .ZN(n5606) );
  NOR4_X1 U817 ( .A1(n5615), .A2(n5616), .A3(n5617), .A4(n5618), .ZN(n5605) );
  OAI221_X1 U818 ( .B1(n2058), .B2(n6082), .C1(n2083), .C2(n6086), .A(n5612), 
        .ZN(n5609) );
  NAND2_X1 U819 ( .A1(n5173), .A2(n5174), .ZN(OUT1[6]) );
  NOR4_X1 U820 ( .A1(n5175), .A2(n5176), .A3(n5177), .A4(n5178), .ZN(n5174) );
  NOR4_X1 U821 ( .A1(n5183), .A2(n5184), .A3(n5185), .A4(n5186), .ZN(n5173) );
  OAI221_X1 U822 ( .B1(n2062), .B2(n6078), .C1(n2090), .C2(n6086), .A(n5180), 
        .ZN(n5177) );
  NAND2_X1 U823 ( .A1(n5389), .A2(n5390), .ZN(OUT1[24]) );
  NOR4_X1 U824 ( .A1(n5391), .A2(n5392), .A3(n5393), .A4(n5394), .ZN(n5390) );
  NOR4_X1 U825 ( .A1(n5399), .A2(n5400), .A3(n5401), .A4(n5402), .ZN(n5389) );
  OAI221_X1 U826 ( .B1(n2047), .B2(n6081), .C1(n2072), .C2(n6089), .A(n5396), 
        .ZN(n5393) );
  NAND2_X1 U827 ( .A1(n5443), .A2(n5444), .ZN(OUT1[21]) );
  NOR4_X1 U828 ( .A1(n5445), .A2(n5446), .A3(n5447), .A4(n5448), .ZN(n5444) );
  NOR4_X1 U829 ( .A1(n5453), .A2(n5454), .A3(n5455), .A4(n5456), .ZN(n5443) );
  OAI221_X1 U830 ( .B1(n2050), .B2(n6079), .C1(n2075), .C2(n6088), .A(n5450), 
        .ZN(n5447) );
  NAND2_X1 U831 ( .A1(n5515), .A2(n5516), .ZN(OUT1[18]) );
  NOR4_X1 U832 ( .A1(n5517), .A2(n5518), .A3(n5519), .A4(n5520), .ZN(n5516) );
  NOR4_X1 U833 ( .A1(n5525), .A2(n5526), .A3(n5527), .A4(n5528), .ZN(n5515) );
  OAI221_X1 U834 ( .B1(n2053), .B2(n6079), .C1(n2078), .C2(n6088), .A(n5522), 
        .ZN(n5519) );
  NAND2_X1 U835 ( .A1(n5587), .A2(n5588), .ZN(OUT1[14]) );
  NOR4_X1 U836 ( .A1(n5589), .A2(n5590), .A3(n5591), .A4(n5592), .ZN(n5588) );
  NOR4_X1 U837 ( .A1(n5597), .A2(n5598), .A3(n5599), .A4(n5600), .ZN(n5587) );
  OAI221_X1 U838 ( .B1(n2057), .B2(n6079), .C1(n2082), .C2(n6088), .A(n5594), 
        .ZN(n5591) );
  NAND2_X1 U839 ( .A1(n5155), .A2(n5156), .ZN(OUT1[7]) );
  NOR4_X1 U840 ( .A1(n5157), .A2(n5158), .A3(n5159), .A4(n5160), .ZN(n5156) );
  NOR4_X1 U841 ( .A1(n5165), .A2(n5166), .A3(n5167), .A4(n5168), .ZN(n5155) );
  OAI221_X1 U842 ( .B1(n2061), .B2(n6078), .C1(n2089), .C2(n6086), .A(n5162), 
        .ZN(n5159) );
  NAND2_X1 U843 ( .A1(n5371), .A2(n5372), .ZN(OUT1[25]) );
  NOR4_X1 U844 ( .A1(n5373), .A2(n5374), .A3(n5375), .A4(n5376), .ZN(n5372) );
  NOR4_X1 U845 ( .A1(n5381), .A2(n5382), .A3(n5383), .A4(n5384), .ZN(n5371) );
  OAI221_X1 U846 ( .B1(n2046), .B2(n6081), .C1(n2071), .C2(n6089), .A(n5378), 
        .ZN(n5375) );
  NAND2_X1 U847 ( .A1(n5087), .A2(n5088), .ZN(OUT1[9]) );
  NOR4_X1 U848 ( .A1(n5089), .A2(n5090), .A3(n5091), .A4(n5092), .ZN(n5088) );
  NOR4_X1 U849 ( .A1(n5113), .A2(n5114), .A3(n5115), .A4(n5116), .ZN(n5087) );
  OAI221_X1 U850 ( .B1(n1923), .B2(n6014), .C1(n1960), .C2(n6022), .A(n5110), 
        .ZN(n5089) );
  NAND2_X1 U851 ( .A1(n5425), .A2(n5426), .ZN(OUT1[22]) );
  NOR4_X1 U852 ( .A1(n5427), .A2(n5428), .A3(n5429), .A4(n5430), .ZN(n5426) );
  NOR4_X1 U853 ( .A1(n5435), .A2(n5436), .A3(n5437), .A4(n5438), .ZN(n5425) );
  OAI221_X1 U854 ( .B1(n2049), .B2(n6080), .C1(n2074), .C2(n6089), .A(n5432), 
        .ZN(n5429) );
  NAND2_X1 U855 ( .A1(n5497), .A2(n5498), .ZN(OUT1[19]) );
  NOR4_X1 U856 ( .A1(n5499), .A2(n5500), .A3(n5501), .A4(n5502), .ZN(n5498) );
  NOR4_X1 U857 ( .A1(n5507), .A2(n5508), .A3(n5509), .A4(n5510), .ZN(n5497) );
  OAI221_X1 U858 ( .B1(n2052), .B2(n6082), .C1(n2077), .C2(n6090), .A(n5504), 
        .ZN(n5501) );
  NAND2_X1 U859 ( .A1(n5569), .A2(n5570), .ZN(OUT1[15]) );
  NOR4_X1 U860 ( .A1(n5571), .A2(n5572), .A3(n5573), .A4(n5574), .ZN(n5570) );
  NOR4_X1 U861 ( .A1(n5579), .A2(n5580), .A3(n5581), .A4(n5582), .ZN(n5569) );
  OAI221_X1 U862 ( .B1(n2056), .B2(n6080), .C1(n2081), .C2(n6089), .A(n5576), 
        .ZN(n5573) );
  NAND2_X1 U863 ( .A1(n5137), .A2(n5138), .ZN(OUT1[8]) );
  NOR4_X1 U864 ( .A1(n5139), .A2(n5140), .A3(n5141), .A4(n5142), .ZN(n5138) );
  NOR4_X1 U865 ( .A1(n5147), .A2(n5148), .A3(n5149), .A4(n5150), .ZN(n5137) );
  OAI221_X1 U866 ( .B1(n2060), .B2(n6078), .C1(n2088), .C2(n6089), .A(n5144), 
        .ZN(n5141) );
  NAND2_X1 U867 ( .A1(n5209), .A2(n5210), .ZN(OUT1[4]) );
  NOR4_X1 U868 ( .A1(n5211), .A2(n5212), .A3(n5213), .A4(n5214), .ZN(n5210) );
  NOR4_X1 U869 ( .A1(n5219), .A2(n5220), .A3(n5221), .A4(n5222), .ZN(n5209) );
  OAI221_X1 U870 ( .B1(n2064), .B2(n6083), .C1(n2092), .C2(n6091), .A(n5216), 
        .ZN(n5213) );
  NAND2_X1 U871 ( .A1(n5407), .A2(n5408), .ZN(OUT1[23]) );
  NOR4_X1 U872 ( .A1(n5409), .A2(n5410), .A3(n5411), .A4(n5412), .ZN(n5408) );
  NOR4_X1 U873 ( .A1(n5417), .A2(n5418), .A3(n5419), .A4(n5420), .ZN(n5407) );
  OAI221_X1 U874 ( .B1(n1897), .B2(n6014), .C1(n1946), .C2(n6025), .A(n5416), 
        .ZN(n5409) );
  NAND2_X1 U875 ( .A1(n5479), .A2(n5480), .ZN(OUT1[1]) );
  NOR4_X1 U876 ( .A1(n5481), .A2(n5482), .A3(n5483), .A4(n5484), .ZN(n5480) );
  NOR4_X1 U877 ( .A1(n5489), .A2(n5490), .A3(n5491), .A4(n5492), .ZN(n5479) );
  OAI221_X1 U878 ( .B1(n2067), .B2(n6078), .C1(n2093), .C2(n6087), .A(n5486), 
        .ZN(n5483) );
  NAND2_X1 U879 ( .A1(n5551), .A2(n5552), .ZN(OUT1[16]) );
  NOR4_X1 U880 ( .A1(n5553), .A2(n5554), .A3(n5555), .A4(n5556), .ZN(n5552) );
  NOR4_X1 U881 ( .A1(n5561), .A2(n5562), .A3(n5563), .A4(n5564), .ZN(n5551) );
  OAI221_X1 U882 ( .B1(n2055), .B2(n6080), .C1(n2080), .C2(n6091), .A(n5558), 
        .ZN(n5555) );
  NAND2_X1 U883 ( .A1(n5623), .A2(n5624), .ZN(OUT1[12]) );
  NOR4_X1 U884 ( .A1(n5625), .A2(n5626), .A3(n5627), .A4(n5628), .ZN(n5624) );
  NOR4_X1 U885 ( .A1(n5633), .A2(n5634), .A3(n5635), .A4(n5636), .ZN(n5623) );
  OAI221_X1 U886 ( .B1(n1919), .B2(n6014), .C1(n1957), .C2(n6022), .A(n5632), 
        .ZN(n5625) );
  NAND2_X1 U887 ( .A1(n5191), .A2(n5192), .ZN(OUT1[5]) );
  NOR4_X1 U888 ( .A1(n5193), .A2(n5194), .A3(n5195), .A4(n5196), .ZN(n5192) );
  NOR4_X1 U889 ( .A1(n5201), .A2(n5202), .A3(n5203), .A4(n5204), .ZN(n5191) );
  OAI221_X1 U890 ( .B1(n2063), .B2(n6081), .C1(n2091), .C2(n6091), .A(n5198), 
        .ZN(n5195) );
  NOR3_X1 U891 ( .A1(n5054), .A2(n5053), .A3(n5075), .ZN(n5080) );
  AND2_X1 U892 ( .A1(n5046), .A2(n5051), .ZN(n6325) );
  AND2_X1 U893 ( .A1(n5046), .A2(n5051), .ZN(n6324) );
  AND2_X1 U894 ( .A1(n5046), .A2(n5045), .ZN(n6345) );
  AND2_X1 U895 ( .A1(n5046), .A2(n5045), .ZN(n6344) );
  AND2_X1 U896 ( .A1(n5044), .A2(n5051), .ZN(n6327) );
  AND2_X1 U897 ( .A1(n5044), .A2(n5051), .ZN(n6326) );
  AND2_X1 U898 ( .A1(n5044), .A2(n5045), .ZN(n6347) );
  AND2_X1 U899 ( .A1(n5044), .A2(n5045), .ZN(n6346) );
  AND2_X1 U900 ( .A1(n5046), .A2(n5051), .ZN(n2364) );
  AND2_X1 U901 ( .A1(n5046), .A2(n5045), .ZN(n2357) );
  AND2_X1 U902 ( .A1(n5044), .A2(n5051), .ZN(n2366) );
  AND2_X1 U903 ( .A1(n5044), .A2(n5045), .ZN(n2359) );
  INV_X1 U904 ( .A(n1944), .ZN(n6628) );
  OAI21_X1 U905 ( .B1(n1941), .B2(n1967), .A(n6735), .ZN(n1944) );
  INV_X1 U906 ( .A(n2345), .ZN(n6367) );
  OAI21_X1 U907 ( .B1(n1970), .B2(n2339), .A(n6735), .ZN(n2345) );
  INV_X1 U908 ( .A(n2338), .ZN(n6385) );
  OAI21_X1 U909 ( .B1(n1942), .B2(n2339), .A(n6735), .ZN(n2338) );
  INV_X1 U910 ( .A(n2155), .ZN(n6511) );
  OAI21_X1 U911 ( .B1(n1970), .B2(n2129), .A(RESET), .ZN(n2155) );
  INV_X1 U912 ( .A(n2100), .ZN(n6529) );
  OAI21_X1 U913 ( .B1(n1942), .B2(n2129), .A(RESET), .ZN(n2100) );
  INV_X1 U914 ( .A(n2096), .ZN(n6547) );
  OAI21_X1 U915 ( .B1(n1970), .B2(n2068), .A(RESET), .ZN(n2096) );
  INV_X1 U916 ( .A(n2039), .ZN(n6565) );
  OAI21_X1 U917 ( .B1(n1942), .B2(n2068), .A(RESET), .ZN(n2039) );
  INV_X1 U918 ( .A(n1969), .ZN(n6619) );
  OAI21_X1 U919 ( .B1(n1941), .B2(n1970), .A(n6735), .ZN(n1969) );
  INV_X1 U920 ( .A(n2035), .ZN(n6583) );
  OAI21_X1 U921 ( .B1(n1970), .B2(n2008), .A(n6735), .ZN(n2035) );
  INV_X1 U922 ( .A(n1978), .ZN(n6601) );
  OAI21_X1 U923 ( .B1(n1942), .B2(n2008), .A(RESET), .ZN(n1978) );
  NAND2_X1 U924 ( .A1(n5047), .A2(n5059), .ZN(n2368) );
  NAND2_X1 U925 ( .A1(n5047), .A2(n5058), .ZN(n2369) );
  NAND2_X1 U926 ( .A1(n5052), .A2(n5059), .ZN(n2375) );
  NAND2_X1 U927 ( .A1(n5052), .A2(n5058), .ZN(n2376) );
  NAND2_X1 U928 ( .A1(n2340), .A2(n2341), .ZN(n1942) );
  OAI221_X1 U929 ( .B1(n2128), .B2(n6333), .C1(n2152), .C2(n6341), .A(n4667), 
        .ZN(n4666) );
  AOI22_X1 U930 ( .A1(n2357), .A2(n4668), .B1(n2359), .B2(n4669), .ZN(n4667)
         );
  OAI221_X1 U931 ( .B1(n2273), .B2(n6217), .C1(n2241), .C2(n6225), .A(n4683), 
        .ZN(n4682) );
  AOI22_X1 U932 ( .A1(n6233), .A2(n4684), .B1(n6241), .B2(n4685), .ZN(n4683)
         );
  OAI221_X1 U933 ( .B1(n2124), .B2(n6335), .C1(n2151), .C2(n6343), .A(n2522), 
        .ZN(n2521) );
  AOI22_X1 U934 ( .A1(n6344), .A2(n2523), .B1(n6346), .B2(n2524), .ZN(n2522)
         );
  OAI221_X1 U935 ( .B1(n2269), .B2(n6219), .C1(n2240), .C2(n6227), .A(n2538), 
        .ZN(n2537) );
  AOI22_X1 U936 ( .A1(n6230), .A2(n2539), .B1(n6238), .B2(n2540), .ZN(n2538)
         );
  OAI221_X1 U937 ( .B1(n2123), .B2(n6329), .C1(n2150), .C2(n6338), .A(n2488), 
        .ZN(n2487) );
  AOI22_X1 U938 ( .A1(n6345), .A2(n2489), .B1(n6347), .B2(n2490), .ZN(n2488)
         );
  OAI221_X1 U939 ( .B1(n2268), .B2(n6213), .C1(n2239), .C2(n6222), .A(n2504), 
        .ZN(n2503) );
  AOI22_X1 U940 ( .A1(n6231), .A2(n2505), .B1(n6239), .B2(n2506), .ZN(n2504)
         );
  OAI221_X1 U941 ( .B1(n2122), .B2(n6329), .C1(n2149), .C2(n6338), .A(n2454), 
        .ZN(n2453) );
  AOI22_X1 U942 ( .A1(n2357), .A2(n2455), .B1(n2359), .B2(n2456), .ZN(n2454)
         );
  OAI221_X1 U943 ( .B1(n2267), .B2(n6213), .C1(n2238), .C2(n6222), .A(n2470), 
        .ZN(n2469) );
  AOI22_X1 U944 ( .A1(n6234), .A2(n2471), .B1(n6240), .B2(n2472), .ZN(n2470)
         );
  OAI221_X1 U945 ( .B1(n2121), .B2(n6335), .C1(n2148), .C2(n6343), .A(n2420), 
        .ZN(n2419) );
  AOI22_X1 U946 ( .A1(n6344), .A2(n2421), .B1(n6346), .B2(n2422), .ZN(n2420)
         );
  OAI221_X1 U947 ( .B1(n2266), .B2(n6219), .C1(n2237), .C2(n6227), .A(n2436), 
        .ZN(n2435) );
  AOI22_X1 U948 ( .A1(n6231), .A2(n2437), .B1(n6239), .B2(n2438), .ZN(n2436)
         );
  OAI221_X1 U949 ( .B1(n2119), .B2(n6330), .C1(n2144), .C2(n6339), .A(n4905), 
        .ZN(n4904) );
  AOI22_X1 U950 ( .A1(n6345), .A2(n4906), .B1(n6347), .B2(n4907), .ZN(n4905)
         );
  OAI221_X1 U951 ( .B1(n2264), .B2(n6214), .C1(n2233), .C2(n6223), .A(n4921), 
        .ZN(n4920) );
  AOI22_X1 U952 ( .A1(n6230), .A2(n4922), .B1(n6238), .B2(n4923), .ZN(n4921)
         );
  OAI221_X1 U953 ( .B1(n2118), .B2(n6331), .C1(n2143), .C2(n6341), .A(n4871), 
        .ZN(n4870) );
  AOI22_X1 U954 ( .A1(n2357), .A2(n4872), .B1(n2359), .B2(n4873), .ZN(n4871)
         );
  OAI221_X1 U955 ( .B1(n2263), .B2(n6215), .C1(n2232), .C2(n6225), .A(n4887), 
        .ZN(n4886) );
  AOI22_X1 U956 ( .A1(n6230), .A2(n4888), .B1(n6238), .B2(n4889), .ZN(n4887)
         );
  OAI221_X1 U957 ( .B1(n2117), .B2(n6332), .C1(n2142), .C2(n6338), .A(n4837), 
        .ZN(n4836) );
  AOI22_X1 U958 ( .A1(n6344), .A2(n4838), .B1(n6346), .B2(n4839), .ZN(n4837)
         );
  OAI221_X1 U959 ( .B1(n2262), .B2(n6216), .C1(n2231), .C2(n6222), .A(n4853), 
        .ZN(n4852) );
  AOI22_X1 U960 ( .A1(n6231), .A2(n4854), .B1(n6239), .B2(n4855), .ZN(n4853)
         );
  OAI221_X1 U961 ( .B1(n2116), .B2(n6332), .C1(n2141), .C2(n6339), .A(n4803), 
        .ZN(n4802) );
  AOI22_X1 U962 ( .A1(n6345), .A2(n4804), .B1(n6347), .B2(n4805), .ZN(n4803)
         );
  OAI221_X1 U963 ( .B1(n2261), .B2(n6216), .C1(n2230), .C2(n6223), .A(n4819), 
        .ZN(n4818) );
  AOI22_X1 U964 ( .A1(n6235), .A2(n4820), .B1(n6240), .B2(n4821), .ZN(n4819)
         );
  OAI221_X1 U965 ( .B1(n2115), .B2(n6330), .C1(n2140), .C2(n6343), .A(n4769), 
        .ZN(n4768) );
  AOI22_X1 U966 ( .A1(n2357), .A2(n4770), .B1(n2359), .B2(n4771), .ZN(n4769)
         );
  OAI221_X1 U967 ( .B1(n2260), .B2(n6214), .C1(n2229), .C2(n6227), .A(n4785), 
        .ZN(n4784) );
  AOI22_X1 U968 ( .A1(n6231), .A2(n4786), .B1(n6240), .B2(n4787), .ZN(n4785)
         );
  OAI221_X1 U969 ( .B1(n2114), .B2(n6335), .C1(n2139), .C2(n6339), .A(n4735), 
        .ZN(n4734) );
  AOI22_X1 U970 ( .A1(n6344), .A2(n4736), .B1(n6346), .B2(n4737), .ZN(n4735)
         );
  OAI221_X1 U971 ( .B1(n2259), .B2(n6219), .C1(n2228), .C2(n6223), .A(n4751), 
        .ZN(n4750) );
  AOI22_X1 U972 ( .A1(n6233), .A2(n4752), .B1(n6241), .B2(n4753), .ZN(n4751)
         );
  OAI221_X1 U973 ( .B1(n2113), .B2(n6331), .C1(n2138), .C2(n6340), .A(n4701), 
        .ZN(n4700) );
  AOI22_X1 U974 ( .A1(n6345), .A2(n4702), .B1(n6347), .B2(n4703), .ZN(n4701)
         );
  OAI221_X1 U975 ( .B1(n2258), .B2(n6215), .C1(n2227), .C2(n6224), .A(n4717), 
        .ZN(n4716) );
  AOI22_X1 U976 ( .A1(n6232), .A2(n4718), .B1(n6241), .B2(n4719), .ZN(n4717)
         );
  OAI221_X1 U977 ( .B1(n2112), .B2(n6330), .C1(n2137), .C2(n6339), .A(n4633), 
        .ZN(n4632) );
  AOI22_X1 U978 ( .A1(n6344), .A2(n4634), .B1(n6346), .B2(n4635), .ZN(n4633)
         );
  OAI221_X1 U979 ( .B1(n2257), .B2(n6214), .C1(n2226), .C2(n6223), .A(n4649), 
        .ZN(n4648) );
  AOI22_X1 U980 ( .A1(n6234), .A2(n4650), .B1(n6242), .B2(n4651), .ZN(n4649)
         );
  OAI221_X1 U981 ( .B1(n2111), .B2(n6331), .C1(n2136), .C2(n6341), .A(n4599), 
        .ZN(n4598) );
  AOI22_X1 U982 ( .A1(n6345), .A2(n4600), .B1(n6347), .B2(n4601), .ZN(n4599)
         );
  OAI221_X1 U983 ( .B1(n2256), .B2(n6215), .C1(n2225), .C2(n6225), .A(n4615), 
        .ZN(n4614) );
  AOI22_X1 U984 ( .A1(n6234), .A2(n4616), .B1(n6242), .B2(n4617), .ZN(n4615)
         );
  OAI221_X1 U985 ( .B1(n2110), .B2(n6331), .C1(n2135), .C2(n6338), .A(n4565), 
        .ZN(n4564) );
  AOI22_X1 U986 ( .A1(n2357), .A2(n4566), .B1(n2359), .B2(n4567), .ZN(n4565)
         );
  OAI221_X1 U987 ( .B1(n2255), .B2(n6215), .C1(n2224), .C2(n6222), .A(n4581), 
        .ZN(n4580) );
  AOI22_X1 U988 ( .A1(n6232), .A2(n4582), .B1(n6241), .B2(n4583), .ZN(n4581)
         );
  OAI221_X1 U989 ( .B1(n2109), .B2(n6332), .C1(n2134), .C2(n6340), .A(n4531), 
        .ZN(n4530) );
  AOI22_X1 U990 ( .A1(n6344), .A2(n4532), .B1(n6346), .B2(n4533), .ZN(n4531)
         );
  OAI221_X1 U991 ( .B1(n2254), .B2(n6216), .C1(n2223), .C2(n6224), .A(n4547), 
        .ZN(n4546) );
  AOI22_X1 U992 ( .A1(n6233), .A2(n4548), .B1(n6243), .B2(n4549), .ZN(n4547)
         );
  OAI221_X1 U993 ( .B1(n2108), .B2(n6329), .C1(n2133), .C2(n6342), .A(n4497), 
        .ZN(n4496) );
  AOI22_X1 U994 ( .A1(n6345), .A2(n4498), .B1(n6347), .B2(n4499), .ZN(n4497)
         );
  OAI221_X1 U995 ( .B1(n2253), .B2(n6213), .C1(n2222), .C2(n6226), .A(n4513), 
        .ZN(n4512) );
  AOI22_X1 U996 ( .A1(n6231), .A2(n4514), .B1(n6242), .B2(n4515), .ZN(n4513)
         );
  OAI221_X1 U997 ( .B1(n2107), .B2(n6334), .C1(n2132), .C2(n6338), .A(n4463), 
        .ZN(n4462) );
  AOI22_X1 U998 ( .A1(n2357), .A2(n4464), .B1(n2359), .B2(n4465), .ZN(n4463)
         );
  OAI221_X1 U999 ( .B1(n2252), .B2(n6218), .C1(n2221), .C2(n6222), .A(n4479), 
        .ZN(n4478) );
  AOI22_X1 U1000 ( .A1(n6234), .A2(n4480), .B1(n6242), .B2(n4481), .ZN(n4479)
         );
  OAI221_X1 U1001 ( .B1(n2067), .B2(n6313), .C1(n2093), .C2(n6321), .A(n4670), 
        .ZN(n4665) );
  AOI22_X1 U1002 ( .A1(n2364), .A2(n4671), .B1(n2366), .B2(n4672), .ZN(n4670)
         );
  OAI221_X1 U1003 ( .B1(n2213), .B2(n6185), .C1(n2181), .C2(n6193), .A(n4686), 
        .ZN(n4681) );
  AOI22_X1 U1004 ( .A1(n6201), .A2(n4687), .B1(n6209), .B2(n4688), .ZN(n4686)
         );
  OAI221_X1 U1005 ( .B1(n2064), .B2(n6314), .C1(n2092), .C2(n6322), .A(n2559), 
        .ZN(n2554) );
  AOI22_X1 U1006 ( .A1(n2364), .A2(n2560), .B1(n2366), .B2(n2561), .ZN(n2559)
         );
  OAI221_X1 U1007 ( .B1(n2063), .B2(n6315), .C1(n2091), .C2(n6323), .A(n2525), 
        .ZN(n2520) );
  AOI22_X1 U1008 ( .A1(n6324), .A2(n2526), .B1(n6326), .B2(n2527), .ZN(n2525)
         );
  OAI221_X1 U1009 ( .B1(n2209), .B2(n6187), .C1(n2180), .C2(n6195), .A(n2541), 
        .ZN(n2536) );
  AOI22_X1 U1010 ( .A1(n6198), .A2(n2542), .B1(n6206), .B2(n2543), .ZN(n2541)
         );
  OAI221_X1 U1011 ( .B1(n2062), .B2(n6309), .C1(n2090), .C2(n6318), .A(n2491), 
        .ZN(n2486) );
  AOI22_X1 U1012 ( .A1(n6325), .A2(n2492), .B1(n6327), .B2(n2493), .ZN(n2491)
         );
  OAI221_X1 U1013 ( .B1(n2208), .B2(n6181), .C1(n2179), .C2(n6190), .A(n2507), 
        .ZN(n2502) );
  AOI22_X1 U1014 ( .A1(n6199), .A2(n2508), .B1(n6207), .B2(n2509), .ZN(n2507)
         );
  OAI221_X1 U1015 ( .B1(n2061), .B2(n6309), .C1(n2089), .C2(n6318), .A(n2457), 
        .ZN(n2452) );
  AOI22_X1 U1016 ( .A1(n2364), .A2(n2458), .B1(n2366), .B2(n2459), .ZN(n2457)
         );
  OAI221_X1 U1017 ( .B1(n2207), .B2(n6181), .C1(n2178), .C2(n6190), .A(n2473), 
        .ZN(n2468) );
  AOI22_X1 U1018 ( .A1(n6202), .A2(n2474), .B1(n6208), .B2(n2475), .ZN(n2473)
         );
  OAI221_X1 U1019 ( .B1(n2060), .B2(n6315), .C1(n2088), .C2(n6323), .A(n2423), 
        .ZN(n2418) );
  AOI22_X1 U1020 ( .A1(n6324), .A2(n2424), .B1(n6326), .B2(n2425), .ZN(n2423)
         );
  OAI221_X1 U1021 ( .B1(n2206), .B2(n6187), .C1(n2177), .C2(n6195), .A(n2439), 
        .ZN(n2434) );
  AOI22_X1 U1022 ( .A1(n6199), .A2(n2440), .B1(n6207), .B2(n2441), .ZN(n2439)
         );
  OAI221_X1 U1023 ( .B1(n2059), .B2(n6311), .C1(n2087), .C2(n6320), .A(n2363), 
        .ZN(n2352) );
  AOI22_X1 U1024 ( .A1(n6325), .A2(n2365), .B1(n6327), .B2(n2367), .ZN(n2363)
         );
  OAI221_X1 U1025 ( .B1(n2058), .B2(n6310), .C1(n2083), .C2(n6319), .A(n4908), 
        .ZN(n4903) );
  AOI22_X1 U1026 ( .A1(n6325), .A2(n4909), .B1(n6327), .B2(n4910), .ZN(n4908)
         );
  OAI221_X1 U1027 ( .B1(n2204), .B2(n6182), .C1(n2173), .C2(n6191), .A(n4924), 
        .ZN(n4919) );
  AOI22_X1 U1028 ( .A1(n6198), .A2(n4925), .B1(n6206), .B2(n4926), .ZN(n4924)
         );
  OAI221_X1 U1029 ( .B1(n2057), .B2(n6311), .C1(n2082), .C2(n6321), .A(n4874), 
        .ZN(n4869) );
  AOI22_X1 U1030 ( .A1(n2364), .A2(n4875), .B1(n2366), .B2(n4876), .ZN(n4874)
         );
  OAI221_X1 U1031 ( .B1(n2203), .B2(n6183), .C1(n2172), .C2(n6193), .A(n4890), 
        .ZN(n4885) );
  AOI22_X1 U1032 ( .A1(n6198), .A2(n4891), .B1(n6206), .B2(n4892), .ZN(n4890)
         );
  OAI221_X1 U1033 ( .B1(n2056), .B2(n6312), .C1(n2081), .C2(n6318), .A(n4840), 
        .ZN(n4835) );
  AOI22_X1 U1034 ( .A1(n6324), .A2(n4841), .B1(n6326), .B2(n4842), .ZN(n4840)
         );
  OAI221_X1 U1035 ( .B1(n2202), .B2(n6184), .C1(n2171), .C2(n6190), .A(n4856), 
        .ZN(n4851) );
  AOI22_X1 U1036 ( .A1(n6199), .A2(n4857), .B1(n6207), .B2(n4858), .ZN(n4856)
         );
  OAI221_X1 U1037 ( .B1(n2055), .B2(n6312), .C1(n2080), .C2(n6319), .A(n4806), 
        .ZN(n4801) );
  AOI22_X1 U1038 ( .A1(n6325), .A2(n4807), .B1(n6327), .B2(n4808), .ZN(n4806)
         );
  OAI221_X1 U1039 ( .B1(n2201), .B2(n6184), .C1(n2170), .C2(n6191), .A(n4822), 
        .ZN(n4817) );
  AOI22_X1 U1040 ( .A1(n6203), .A2(n4823), .B1(n6208), .B2(n4824), .ZN(n4822)
         );
  OAI221_X1 U1041 ( .B1(n2054), .B2(n6310), .C1(n2079), .C2(n6323), .A(n4772), 
        .ZN(n4767) );
  AOI22_X1 U1042 ( .A1(n2364), .A2(n4773), .B1(n2366), .B2(n4774), .ZN(n4772)
         );
  OAI221_X1 U1043 ( .B1(n2200), .B2(n6182), .C1(n2169), .C2(n6195), .A(n4788), 
        .ZN(n4783) );
  AOI22_X1 U1044 ( .A1(n6199), .A2(n4789), .B1(n6208), .B2(n4790), .ZN(n4788)
         );
  OAI221_X1 U1045 ( .B1(n2053), .B2(n6315), .C1(n2078), .C2(n6319), .A(n4738), 
        .ZN(n4733) );
  AOI22_X1 U1046 ( .A1(n6324), .A2(n4739), .B1(n6326), .B2(n4740), .ZN(n4738)
         );
  OAI221_X1 U1047 ( .B1(n2199), .B2(n6187), .C1(n2168), .C2(n6191), .A(n4754), 
        .ZN(n4749) );
  AOI22_X1 U1048 ( .A1(n6201), .A2(n4755), .B1(n6209), .B2(n4756), .ZN(n4754)
         );
  OAI221_X1 U1049 ( .B1(n2052), .B2(n6313), .C1(n2077), .C2(n6320), .A(n4704), 
        .ZN(n4699) );
  AOI22_X1 U1050 ( .A1(n6325), .A2(n4705), .B1(n6327), .B2(n4706), .ZN(n4704)
         );
  OAI221_X1 U1051 ( .B1(n2198), .B2(n6183), .C1(n2167), .C2(n6192), .A(n4720), 
        .ZN(n4715) );
  AOI22_X1 U1052 ( .A1(n6200), .A2(n4721), .B1(n6209), .B2(n4722), .ZN(n4720)
         );
  OAI221_X1 U1053 ( .B1(n2051), .B2(n6310), .C1(n2076), .C2(n6319), .A(n4636), 
        .ZN(n4631) );
  AOI22_X1 U1054 ( .A1(n6324), .A2(n4637), .B1(n6326), .B2(n4638), .ZN(n4636)
         );
  OAI221_X1 U1055 ( .B1(n2197), .B2(n6182), .C1(n2166), .C2(n6191), .A(n4652), 
        .ZN(n4647) );
  AOI22_X1 U1056 ( .A1(n6202), .A2(n4653), .B1(n6210), .B2(n4654), .ZN(n4652)
         );
  OAI221_X1 U1057 ( .B1(n2050), .B2(n6311), .C1(n2075), .C2(n6321), .A(n4602), 
        .ZN(n4597) );
  AOI22_X1 U1058 ( .A1(n6325), .A2(n4603), .B1(n6327), .B2(n4604), .ZN(n4602)
         );
  OAI221_X1 U1059 ( .B1(n2196), .B2(n6183), .C1(n2165), .C2(n6193), .A(n4618), 
        .ZN(n4613) );
  AOI22_X1 U1060 ( .A1(n6202), .A2(n4619), .B1(n6210), .B2(n4620), .ZN(n4618)
         );
  OAI221_X1 U1061 ( .B1(n2049), .B2(n6311), .C1(n2074), .C2(n6318), .A(n4568), 
        .ZN(n4563) );
  AOI22_X1 U1062 ( .A1(n2364), .A2(n4569), .B1(n2366), .B2(n4570), .ZN(n4568)
         );
  OAI221_X1 U1063 ( .B1(n2195), .B2(n6183), .C1(n2164), .C2(n6190), .A(n4584), 
        .ZN(n4579) );
  AOI22_X1 U1064 ( .A1(n6200), .A2(n4585), .B1(n6209), .B2(n4586), .ZN(n4584)
         );
  OAI221_X1 U1065 ( .B1(n2048), .B2(n6312), .C1(n2073), .C2(n6320), .A(n4534), 
        .ZN(n4529) );
  AOI22_X1 U1066 ( .A1(n6324), .A2(n4535), .B1(n6326), .B2(n4536), .ZN(n4534)
         );
  OAI221_X1 U1067 ( .B1(n2194), .B2(n6184), .C1(n2163), .C2(n6192), .A(n4550), 
        .ZN(n4545) );
  AOI22_X1 U1068 ( .A1(n6201), .A2(n4551), .B1(n6211), .B2(n4552), .ZN(n4550)
         );
  OAI221_X1 U1069 ( .B1(n2047), .B2(n6309), .C1(n2072), .C2(n6322), .A(n4500), 
        .ZN(n4495) );
  AOI22_X1 U1070 ( .A1(n6325), .A2(n4501), .B1(n6327), .B2(n4502), .ZN(n4500)
         );
  OAI221_X1 U1071 ( .B1(n2193), .B2(n6181), .C1(n2162), .C2(n6194), .A(n4516), 
        .ZN(n4511) );
  AOI22_X1 U1072 ( .A1(n6199), .A2(n4517), .B1(n6210), .B2(n4518), .ZN(n4516)
         );
  OAI221_X1 U1073 ( .B1(n2046), .B2(n6313), .C1(n2071), .C2(n6318), .A(n4466), 
        .ZN(n4461) );
  AOI22_X1 U1074 ( .A1(n2364), .A2(n4467), .B1(n2366), .B2(n4468), .ZN(n4466)
         );
  OAI221_X1 U1075 ( .B1(n2192), .B2(n6186), .C1(n2161), .C2(n6190), .A(n4482), 
        .ZN(n4477) );
  AOI22_X1 U1076 ( .A1(n6202), .A2(n4483), .B1(n6210), .B2(n4484), .ZN(n4482)
         );
  OAI221_X1 U1077 ( .B1(n2007), .B2(n6280), .C1(n2032), .C2(n6289), .A(n4673), 
        .ZN(n4664) );
  AOI22_X1 U1078 ( .A1(n6293), .A2(n4674), .B1(n6305), .B2(n4675), .ZN(n4673)
         );
  OAI221_X1 U1079 ( .B1(n2307), .B2(n6153), .C1(n2331), .C2(n6161), .A(n4689), 
        .ZN(n4680) );
  AOI22_X1 U1080 ( .A1(n6169), .A2(n4690), .B1(n6177), .B2(n4691), .ZN(n4689)
         );
  OAI221_X1 U1081 ( .B1(n2004), .B2(n6282), .C1(n2031), .C2(n6290), .A(n2562), 
        .ZN(n2553) );
  AOI22_X1 U1082 ( .A1(n6294), .A2(n2563), .B1(n6301), .B2(n2564), .ZN(n2562)
         );
  OAI221_X1 U1083 ( .B1(n2003), .B2(n6283), .C1(n2030), .C2(n6291), .A(n2528), 
        .ZN(n2519) );
  AOI22_X1 U1084 ( .A1(n6295), .A2(n2529), .B1(n6302), .B2(n2530), .ZN(n2528)
         );
  OAI221_X1 U1085 ( .B1(n2303), .B2(n6155), .C1(n2330), .C2(n6163), .A(n2544), 
        .ZN(n2535) );
  AOI22_X1 U1086 ( .A1(n6166), .A2(n2545), .B1(n6174), .B2(n2546), .ZN(n2544)
         );
  OAI221_X1 U1087 ( .B1(n2002), .B2(n6278), .C1(n2029), .C2(n6285), .A(n2494), 
        .ZN(n2485) );
  AOI22_X1 U1088 ( .A1(n6296), .A2(n2495), .B1(n6303), .B2(n2496), .ZN(n2494)
         );
  OAI221_X1 U1089 ( .B1(n2302), .B2(n6149), .C1(n2329), .C2(n6158), .A(n2510), 
        .ZN(n2501) );
  AOI22_X1 U1090 ( .A1(n6167), .A2(n2511), .B1(n6175), .B2(n2512), .ZN(n2510)
         );
  OAI221_X1 U1091 ( .B1(n2001), .B2(n6283), .C1(n2028), .C2(n6291), .A(n2460), 
        .ZN(n2451) );
  AOI22_X1 U1092 ( .A1(n6297), .A2(n2461), .B1(n6304), .B2(n2462), .ZN(n2460)
         );
  OAI221_X1 U1093 ( .B1(n2301), .B2(n6149), .C1(n2328), .C2(n6158), .A(n2476), 
        .ZN(n2467) );
  AOI22_X1 U1094 ( .A1(n6170), .A2(n2477), .B1(n6176), .B2(n2478), .ZN(n2476)
         );
  OAI221_X1 U1095 ( .B1(n2300), .B2(n6155), .C1(n2327), .C2(n6163), .A(n2442), 
        .ZN(n2433) );
  AOI22_X1 U1096 ( .A1(n6167), .A2(n2443), .B1(n6175), .B2(n2444), .ZN(n2442)
         );
  OAI221_X1 U1097 ( .B1(n1999), .B2(n6279), .C1(n2027), .C2(n6285), .A(n2370), 
        .ZN(n2351) );
  AOI22_X1 U1098 ( .A1(n6298), .A2(n2372), .B1(n6305), .B2(n2374), .ZN(n2370)
         );
  OAI221_X1 U1099 ( .B1(n1998), .B2(n6279), .C1(n2024), .C2(n6285), .A(n4945), 
        .ZN(n4936) );
  AOI22_X1 U1100 ( .A1(n6295), .A2(n4946), .B1(n6302), .B2(n4947), .ZN(n4945)
         );
  OAI221_X1 U1101 ( .B1(n1997), .B2(n6278), .C1(n2023), .C2(n6286), .A(n4911), 
        .ZN(n4902) );
  AOI22_X1 U1102 ( .A1(n6294), .A2(n4912), .B1(n6301), .B2(n4913), .ZN(n4911)
         );
  OAI221_X1 U1103 ( .B1(n2298), .B2(n6150), .C1(n2323), .C2(n6159), .A(n4927), 
        .ZN(n4918) );
  AOI22_X1 U1104 ( .A1(n6166), .A2(n4928), .B1(n6174), .B2(n4929), .ZN(n4927)
         );
  OAI221_X1 U1105 ( .B1(n1996), .B2(n6281), .C1(n2022), .C2(n6287), .A(n4877), 
        .ZN(n4868) );
  AOI22_X1 U1106 ( .A1(n6295), .A2(n4878), .B1(n6302), .B2(n4879), .ZN(n4877)
         );
  OAI221_X1 U1107 ( .B1(n2297), .B2(n6151), .C1(n2322), .C2(n6161), .A(n4893), 
        .ZN(n4884) );
  AOI22_X1 U1108 ( .A1(n6166), .A2(n4894), .B1(n6174), .B2(n4895), .ZN(n4893)
         );
  OAI221_X1 U1109 ( .B1(n1995), .B2(n6279), .C1(n2021), .C2(n6287), .A(n4843), 
        .ZN(n4834) );
  AOI22_X1 U1110 ( .A1(n6296), .A2(n4844), .B1(n6303), .B2(n4845), .ZN(n4843)
         );
  OAI221_X1 U1111 ( .B1(n2296), .B2(n6152), .C1(n2321), .C2(n6158), .A(n4859), 
        .ZN(n4850) );
  AOI22_X1 U1112 ( .A1(n6167), .A2(n4860), .B1(n6175), .B2(n4861), .ZN(n4859)
         );
  OAI221_X1 U1113 ( .B1(n1994), .B2(n6278), .C1(n2020), .C2(n6287), .A(n4809), 
        .ZN(n4800) );
  AOI22_X1 U1114 ( .A1(n6297), .A2(n4810), .B1(n6304), .B2(n4811), .ZN(n4809)
         );
  OAI221_X1 U1115 ( .B1(n2295), .B2(n6152), .C1(n2320), .C2(n6159), .A(n4825), 
        .ZN(n4816) );
  AOI22_X1 U1116 ( .A1(n6171), .A2(n4826), .B1(n6176), .B2(n4827), .ZN(n4825)
         );
  OAI221_X1 U1117 ( .B1(n1993), .B2(n6278), .C1(n2019), .C2(n6291), .A(n4775), 
        .ZN(n4766) );
  AOI22_X1 U1118 ( .A1(n6297), .A2(n4776), .B1(n6304), .B2(n4777), .ZN(n4775)
         );
  OAI221_X1 U1119 ( .B1(n2294), .B2(n6150), .C1(n2319), .C2(n6163), .A(n4791), 
        .ZN(n4782) );
  AOI22_X1 U1120 ( .A1(n6167), .A2(n4792), .B1(n6176), .B2(n4793), .ZN(n4791)
         );
  OAI221_X1 U1121 ( .B1(n1992), .B2(n6282), .C1(n2018), .C2(n6286), .A(n4741), 
        .ZN(n4732) );
  AOI22_X1 U1122 ( .A1(n6298), .A2(n4742), .B1(n6305), .B2(n4743), .ZN(n4741)
         );
  OAI221_X1 U1123 ( .B1(n2293), .B2(n6155), .C1(n2318), .C2(n6159), .A(n4757), 
        .ZN(n4748) );
  AOI22_X1 U1124 ( .A1(n6169), .A2(n4758), .B1(n6177), .B2(n4759), .ZN(n4757)
         );
  OAI221_X1 U1125 ( .B1(n1991), .B2(n6280), .C1(n2017), .C2(n6288), .A(n4707), 
        .ZN(n4698) );
  AOI22_X1 U1126 ( .A1(n6298), .A2(n4708), .B1(n6307), .B2(n4709), .ZN(n4707)
         );
  OAI221_X1 U1127 ( .B1(n2292), .B2(n6151), .C1(n2317), .C2(n6160), .A(n4723), 
        .ZN(n4714) );
  AOI22_X1 U1128 ( .A1(n6168), .A2(n4724), .B1(n6177), .B2(n4725), .ZN(n4723)
         );
  OAI221_X1 U1129 ( .B1(n1990), .B2(n6279), .C1(n2016), .C2(n6286), .A(n4639), 
        .ZN(n4630) );
  AOI22_X1 U1130 ( .A1(n6299), .A2(n4640), .B1(n6306), .B2(n4641), .ZN(n4639)
         );
  OAI221_X1 U1131 ( .B1(n2291), .B2(n6150), .C1(n2316), .C2(n6159), .A(n4655), 
        .ZN(n4646) );
  AOI22_X1 U1132 ( .A1(n6170), .A2(n4656), .B1(n6178), .B2(n4657), .ZN(n4655)
         );
  OAI221_X1 U1133 ( .B1(n1989), .B2(n6281), .C1(n2015), .C2(n6287), .A(n4605), 
        .ZN(n4596) );
  AOI22_X1 U1134 ( .A1(n6299), .A2(n4606), .B1(n6306), .B2(n4607), .ZN(n4605)
         );
  OAI221_X1 U1135 ( .B1(n2290), .B2(n6151), .C1(n2315), .C2(n6161), .A(n4621), 
        .ZN(n4612) );
  AOI22_X1 U1136 ( .A1(n6170), .A2(n4622), .B1(n6178), .B2(n4623), .ZN(n4621)
         );
  OAI221_X1 U1137 ( .B1(n1988), .B2(n6280), .C1(n2014), .C2(n6287), .A(n4571), 
        .ZN(n4562) );
  AOI22_X1 U1138 ( .A1(n6298), .A2(n4572), .B1(n6305), .B2(n4573), .ZN(n4571)
         );
  OAI221_X1 U1139 ( .B1(n2289), .B2(n6151), .C1(n2314), .C2(n6158), .A(n4587), 
        .ZN(n4578) );
  AOI22_X1 U1140 ( .A1(n6168), .A2(n4588), .B1(n6177), .B2(n4589), .ZN(n4587)
         );
  OAI221_X1 U1141 ( .B1(n1987), .B2(n6278), .C1(n2013), .C2(n6287), .A(n4537), 
        .ZN(n4528) );
  AOI22_X1 U1142 ( .A1(n6294), .A2(n4538), .B1(n6305), .B2(n4539), .ZN(n4537)
         );
  OAI221_X1 U1143 ( .B1(n2288), .B2(n6152), .C1(n2313), .C2(n6160), .A(n4553), 
        .ZN(n4544) );
  AOI22_X1 U1144 ( .A1(n6169), .A2(n4554), .B1(n6179), .B2(n4555), .ZN(n4553)
         );
  OAI221_X1 U1145 ( .B1(n1986), .B2(n6279), .C1(n2012), .C2(n6290), .A(n4503), 
        .ZN(n4494) );
  AOI22_X1 U1146 ( .A1(n6295), .A2(n4504), .B1(n6306), .B2(n4505), .ZN(n4503)
         );
  OAI221_X1 U1147 ( .B1(n2287), .B2(n6149), .C1(n2312), .C2(n6162), .A(n4519), 
        .ZN(n4510) );
  AOI22_X1 U1148 ( .A1(n6167), .A2(n4520), .B1(n6178), .B2(n4521), .ZN(n4519)
         );
  OAI221_X1 U1149 ( .B1(n1985), .B2(n6283), .C1(n2011), .C2(n6285), .A(n4469), 
        .ZN(n4460) );
  AOI22_X1 U1150 ( .A1(n6299), .A2(n4470), .B1(n6306), .B2(n4471), .ZN(n4469)
         );
  OAI221_X1 U1151 ( .B1(n2286), .B2(n6154), .C1(n2311), .C2(n6158), .A(n4485), 
        .ZN(n4476) );
  AOI22_X1 U1152 ( .A1(n6170), .A2(n4486), .B1(n6178), .B2(n4487), .ZN(n4485)
         );
  OAI221_X1 U1153 ( .B1(n1939), .B2(n6248), .C1(n1965), .C2(n6257), .A(n4676), 
        .ZN(n4663) );
  AOI22_X1 U1154 ( .A1(n6265), .A2(n4677), .B1(n6273), .B2(n4678), .ZN(n4676)
         );
  OAI221_X1 U1155 ( .B1(n1933), .B2(n6250), .C1(n1964), .C2(n6258), .A(n2565), 
        .ZN(n2552) );
  AOI22_X1 U1156 ( .A1(n6262), .A2(n2566), .B1(n6269), .B2(n2567), .ZN(n2565)
         );
  OAI221_X1 U1157 ( .B1(n1931), .B2(n6251), .C1(n1963), .C2(n6259), .A(n2531), 
        .ZN(n2518) );
  AOI22_X1 U1158 ( .A1(n6262), .A2(n2532), .B1(n6270), .B2(n2533), .ZN(n2531)
         );
  OAI221_X1 U1159 ( .B1(n1929), .B2(n6246), .C1(n1962), .C2(n6253), .A(n2497), 
        .ZN(n2484) );
  AOI22_X1 U1160 ( .A1(n6263), .A2(n2498), .B1(n6271), .B2(n2499), .ZN(n2497)
         );
  OAI221_X1 U1161 ( .B1(n1927), .B2(n6250), .C1(n1961), .C2(n6258), .A(n2463), 
        .ZN(n2450) );
  AOI22_X1 U1162 ( .A1(n6264), .A2(n2464), .B1(n6272), .B2(n2465), .ZN(n2463)
         );
  OAI221_X1 U1163 ( .B1(n1923), .B2(n6246), .C1(n1960), .C2(n6253), .A(n2377), 
        .ZN(n2350) );
  AOI22_X1 U1164 ( .A1(n6265), .A2(n2379), .B1(n6273), .B2(n2381), .ZN(n2377)
         );
  OAI221_X1 U1165 ( .B1(n1919), .B2(n6246), .C1(n1957), .C2(n6253), .A(n4948), 
        .ZN(n4935) );
  AOI22_X1 U1166 ( .A1(n6262), .A2(n4949), .B1(n6270), .B2(n4950), .ZN(n4948)
         );
  OAI221_X1 U1167 ( .B1(n1917), .B2(n6247), .C1(n1956), .C2(n6253), .A(n4914), 
        .ZN(n4901) );
  AOI22_X1 U1168 ( .A1(n6262), .A2(n4915), .B1(n6269), .B2(n4916), .ZN(n4914)
         );
  OAI221_X1 U1169 ( .B1(n1915), .B2(n6249), .C1(n1955), .C2(n6254), .A(n4880), 
        .ZN(n4867) );
  AOI22_X1 U1170 ( .A1(n6266), .A2(n4881), .B1(n6270), .B2(n4882), .ZN(n4880)
         );
  OAI221_X1 U1171 ( .B1(n1913), .B2(n6247), .C1(n1954), .C2(n6255), .A(n4846), 
        .ZN(n4833) );
  AOI22_X1 U1172 ( .A1(n6263), .A2(n4847), .B1(n6271), .B2(n4848), .ZN(n4846)
         );
  OAI221_X1 U1173 ( .B1(n1911), .B2(n6246), .C1(n1953), .C2(n6255), .A(n4812), 
        .ZN(n4799) );
  AOI22_X1 U1174 ( .A1(n6264), .A2(n4813), .B1(n6272), .B2(n4814), .ZN(n4812)
         );
  OAI221_X1 U1175 ( .B1(n1909), .B2(n6250), .C1(n1952), .C2(n6256), .A(n4778), 
        .ZN(n4765) );
  AOI22_X1 U1176 ( .A1(n6264), .A2(n4779), .B1(n6271), .B2(n4780), .ZN(n4778)
         );
  OAI221_X1 U1177 ( .B1(n1907), .B2(n6247), .C1(n1951), .C2(n6257), .A(n4744), 
        .ZN(n4731) );
  AOI22_X1 U1178 ( .A1(n6265), .A2(n4745), .B1(n6273), .B2(n4746), .ZN(n4744)
         );
  OAI221_X1 U1179 ( .B1(n1905), .B2(n6248), .C1(n1950), .C2(n6256), .A(n4710), 
        .ZN(n4697) );
  AOI22_X1 U1180 ( .A1(n6261), .A2(n4711), .B1(n6273), .B2(n4712), .ZN(n4710)
         );
  OAI221_X1 U1181 ( .B1(n1903), .B2(n6247), .C1(n1949), .C2(n6253), .A(n4642), 
        .ZN(n4629) );
  AOI22_X1 U1182 ( .A1(n6266), .A2(n4643), .B1(n6274), .B2(n4644), .ZN(n4642)
         );
  OAI221_X1 U1183 ( .B1(n1901), .B2(n6249), .C1(n1948), .C2(n6254), .A(n4608), 
        .ZN(n4595) );
  AOI22_X1 U1184 ( .A1(n6266), .A2(n4609), .B1(n6274), .B2(n4610), .ZN(n4608)
         );
  OAI221_X1 U1185 ( .B1(n1899), .B2(n6247), .C1(n1947), .C2(n6255), .A(n4574), 
        .ZN(n4561) );
  AOI22_X1 U1186 ( .A1(n6261), .A2(n4575), .B1(n6275), .B2(n4576), .ZN(n4574)
         );
  OAI221_X1 U1187 ( .B1(n1897), .B2(n6248), .C1(n1946), .C2(n6254), .A(n4540), 
        .ZN(n4527) );
  AOI22_X1 U1188 ( .A1(n6265), .A2(n4541), .B1(n6273), .B2(n4542), .ZN(n4540)
         );
  OAI221_X1 U1189 ( .B1(n1895), .B2(n6251), .C1(n1945), .C2(n6259), .A(n4506), 
        .ZN(n4493) );
  AOI22_X1 U1190 ( .A1(n6266), .A2(n4507), .B1(n6274), .B2(n4508), .ZN(n4506)
         );
  NAND2_X1 U1191 ( .A1(n5046), .A2(n5047), .ZN(n2354) );
  NAND2_X1 U1192 ( .A1(n5044), .A2(n5047), .ZN(n2355) );
  NAND2_X1 U1193 ( .A1(n5046), .A2(n5052), .ZN(n2361) );
  NAND2_X1 U1194 ( .A1(n5044), .A2(n5052), .ZN(n2362) );
  NAND2_X1 U1195 ( .A1(n5071), .A2(n5047), .ZN(n2386) );
  NAND2_X1 U1196 ( .A1(n5070), .A2(n5047), .ZN(n2387) );
  NAND2_X1 U1197 ( .A1(n5080), .A2(n5047), .ZN(n2407) );
  NAND2_X1 U1198 ( .A1(n5079), .A2(n5047), .ZN(n2408) );
  NAND2_X1 U1199 ( .A1(n5071), .A2(n5052), .ZN(n2393) );
  NAND2_X1 U1200 ( .A1(n5070), .A2(n5052), .ZN(n2394) );
  NAND2_X1 U1201 ( .A1(n5079), .A2(n5052), .ZN(n2400) );
  NAND2_X1 U1202 ( .A1(n5080), .A2(n5052), .ZN(n2401) );
  OAI22_X1 U1203 ( .A1(n6406), .A2(n6646), .B1(n6404), .B2(n2330), .ZN(n2854)
         );
  OAI22_X1 U1204 ( .A1(n6406), .A2(n6649), .B1(n2310), .B2(n2329), .ZN(n2855)
         );
  OAI22_X1 U1205 ( .A1(n6406), .A2(n6652), .B1(n6404), .B2(n2328), .ZN(n2856)
         );
  OAI22_X1 U1206 ( .A1(n6406), .A2(n6655), .B1(n2310), .B2(n2327), .ZN(n2857)
         );
  OAI22_X1 U1207 ( .A1(n6407), .A2(n6661), .B1(n6404), .B2(n2326), .ZN(n2859)
         );
  OAI22_X1 U1208 ( .A1(n6407), .A2(n6664), .B1(n2310), .B2(n2325), .ZN(n2860)
         );
  OAI22_X1 U1209 ( .A1(n6407), .A2(n6667), .B1(n2310), .B2(n2324), .ZN(n2861)
         );
  OAI22_X1 U1210 ( .A1(n6414), .A2(n6637), .B1(n6413), .B2(n2306), .ZN(n2883)
         );
  OAI22_X1 U1211 ( .A1(n6414), .A2(n6640), .B1(n2279), .B2(n2305), .ZN(n2884)
         );
  OAI22_X1 U1212 ( .A1(n6414), .A2(n6643), .B1(n6413), .B2(n2304), .ZN(n2885)
         );
  OAI22_X1 U1213 ( .A1(n6415), .A2(n6646), .B1(n2279), .B2(n2303), .ZN(n2886)
         );
  OAI22_X1 U1214 ( .A1(n6415), .A2(n6649), .B1(n6413), .B2(n2302), .ZN(n2887)
         );
  OAI22_X1 U1215 ( .A1(n6415), .A2(n6652), .B1(n2279), .B2(n2301), .ZN(n2888)
         );
  OAI22_X1 U1216 ( .A1(n6415), .A2(n6655), .B1(n2279), .B2(n2300), .ZN(n2889)
         );
  OAI22_X1 U1217 ( .A1(n6441), .A2(n6636), .B1(n6440), .B2(n2272), .ZN(n2979)
         );
  OAI22_X1 U1218 ( .A1(n6441), .A2(n6639), .B1(n2245), .B2(n2271), .ZN(n2980)
         );
  OAI22_X1 U1219 ( .A1(n6441), .A2(n6642), .B1(n6440), .B2(n2270), .ZN(n2981)
         );
  OAI22_X1 U1220 ( .A1(n6442), .A2(n6645), .B1(n2245), .B2(n2269), .ZN(n2982)
         );
  OAI22_X1 U1221 ( .A1(n6442), .A2(n6648), .B1(n6440), .B2(n2268), .ZN(n2983)
         );
  OAI22_X1 U1222 ( .A1(n6442), .A2(n6651), .B1(n2245), .B2(n2267), .ZN(n2984)
         );
  OAI22_X1 U1223 ( .A1(n6442), .A2(n6654), .B1(n2245), .B2(n2266), .ZN(n2985)
         );
  OAI22_X1 U1224 ( .A1(n6451), .A2(n6645), .B1(n6449), .B2(n2240), .ZN(n3014)
         );
  OAI22_X1 U1225 ( .A1(n6451), .A2(n6648), .B1(n2220), .B2(n2239), .ZN(n3015)
         );
  OAI22_X1 U1226 ( .A1(n6451), .A2(n6651), .B1(n6449), .B2(n2238), .ZN(n3016)
         );
  OAI22_X1 U1227 ( .A1(n6451), .A2(n6654), .B1(n2220), .B2(n2237), .ZN(n3017)
         );
  OAI22_X1 U1228 ( .A1(n6452), .A2(n6660), .B1(n6449), .B2(n2236), .ZN(n3019)
         );
  OAI22_X1 U1229 ( .A1(n6452), .A2(n6663), .B1(n2220), .B2(n2235), .ZN(n3020)
         );
  OAI22_X1 U1230 ( .A1(n6452), .A2(n6666), .B1(n2220), .B2(n2234), .ZN(n3021)
         );
  OAI22_X1 U1231 ( .A1(n6477), .A2(n6636), .B1(n6476), .B2(n2212), .ZN(n3107)
         );
  OAI22_X1 U1232 ( .A1(n6477), .A2(n6639), .B1(n2185), .B2(n2211), .ZN(n3108)
         );
  OAI22_X1 U1233 ( .A1(n6477), .A2(n6642), .B1(n6476), .B2(n2210), .ZN(n3109)
         );
  OAI22_X1 U1234 ( .A1(n6478), .A2(n6645), .B1(n2185), .B2(n2209), .ZN(n3110)
         );
  OAI22_X1 U1235 ( .A1(n6478), .A2(n6648), .B1(n6476), .B2(n2208), .ZN(n3111)
         );
  OAI22_X1 U1236 ( .A1(n6478), .A2(n6651), .B1(n2185), .B2(n2207), .ZN(n3112)
         );
  OAI22_X1 U1237 ( .A1(n6478), .A2(n6654), .B1(n2185), .B2(n2206), .ZN(n3113)
         );
  OAI22_X1 U1238 ( .A1(n6487), .A2(n6645), .B1(n6485), .B2(n2180), .ZN(n3142)
         );
  OAI22_X1 U1239 ( .A1(n6487), .A2(n6648), .B1(n2160), .B2(n2179), .ZN(n3143)
         );
  OAI22_X1 U1240 ( .A1(n6487), .A2(n6651), .B1(n6485), .B2(n2178), .ZN(n3144)
         );
  OAI22_X1 U1241 ( .A1(n6487), .A2(n6654), .B1(n2160), .B2(n2177), .ZN(n3145)
         );
  OAI22_X1 U1242 ( .A1(n6488), .A2(n6660), .B1(n6485), .B2(n2176), .ZN(n3147)
         );
  OAI22_X1 U1243 ( .A1(n6488), .A2(n6663), .B1(n2160), .B2(n2175), .ZN(n3148)
         );
  OAI22_X1 U1244 ( .A1(n6488), .A2(n6666), .B1(n2160), .B2(n2174), .ZN(n3149)
         );
  OAI22_X1 U1245 ( .A1(n6514), .A2(n6645), .B1(n6512), .B2(n2151), .ZN(n3238)
         );
  OAI22_X1 U1246 ( .A1(n6514), .A2(n6648), .B1(n2131), .B2(n2150), .ZN(n3239)
         );
  OAI22_X1 U1247 ( .A1(n6514), .A2(n6651), .B1(n6512), .B2(n2149), .ZN(n3240)
         );
  OAI22_X1 U1248 ( .A1(n6514), .A2(n6654), .B1(n2131), .B2(n2148), .ZN(n3241)
         );
  OAI22_X1 U1249 ( .A1(n6515), .A2(n6660), .B1(n6512), .B2(n2147), .ZN(n3243)
         );
  OAI22_X1 U1250 ( .A1(n6515), .A2(n6663), .B1(n2131), .B2(n2146), .ZN(n3244)
         );
  OAI22_X1 U1251 ( .A1(n6515), .A2(n6666), .B1(n2131), .B2(n2145), .ZN(n3245)
         );
  OAI22_X1 U1252 ( .A1(n6522), .A2(n6636), .B1(n6521), .B2(n2127), .ZN(n3267)
         );
  OAI22_X1 U1253 ( .A1(n6522), .A2(n6639), .B1(n2100), .B2(n2126), .ZN(n3268)
         );
  OAI22_X1 U1254 ( .A1(n6522), .A2(n6642), .B1(n6521), .B2(n2125), .ZN(n3269)
         );
  OAI22_X1 U1255 ( .A1(n6523), .A2(n6645), .B1(n2100), .B2(n2124), .ZN(n3270)
         );
  OAI22_X1 U1256 ( .A1(n6523), .A2(n6648), .B1(n6521), .B2(n2123), .ZN(n3271)
         );
  OAI22_X1 U1257 ( .A1(n6523), .A2(n6651), .B1(n2100), .B2(n2122), .ZN(n3272)
         );
  OAI22_X1 U1258 ( .A1(n6523), .A2(n6654), .B1(n2100), .B2(n2121), .ZN(n3273)
         );
  OAI22_X1 U1259 ( .A1(n6549), .A2(n6641), .B1(n6548), .B2(n2092), .ZN(n3365)
         );
  OAI22_X1 U1260 ( .A1(n6550), .A2(n6644), .B1(n2070), .B2(n2091), .ZN(n3366)
         );
  OAI22_X1 U1261 ( .A1(n6550), .A2(n6647), .B1(n6548), .B2(n2090), .ZN(n3367)
         );
  OAI22_X1 U1262 ( .A1(n6550), .A2(n6650), .B1(n2070), .B2(n2089), .ZN(n3368)
         );
  OAI22_X1 U1263 ( .A1(n6550), .A2(n6653), .B1(n6548), .B2(n2088), .ZN(n3369)
         );
  OAI22_X1 U1264 ( .A1(n6550), .A2(n6656), .B1(n2070), .B2(n2087), .ZN(n3370)
         );
  OAI22_X1 U1265 ( .A1(n6551), .A2(n6659), .B1(n2070), .B2(n2086), .ZN(n3371)
         );
  OAI22_X1 U1266 ( .A1(n6558), .A2(n6635), .B1(n6557), .B2(n2066), .ZN(n3395)
         );
  OAI22_X1 U1267 ( .A1(n6558), .A2(n6638), .B1(n2039), .B2(n2065), .ZN(n3396)
         );
  OAI22_X1 U1268 ( .A1(n6558), .A2(n6641), .B1(n6557), .B2(n2064), .ZN(n3397)
         );
  OAI22_X1 U1269 ( .A1(n6559), .A2(n6644), .B1(n2039), .B2(n2063), .ZN(n3398)
         );
  OAI22_X1 U1270 ( .A1(n6559), .A2(n6647), .B1(n6557), .B2(n2062), .ZN(n3399)
         );
  OAI22_X1 U1271 ( .A1(n6559), .A2(n6650), .B1(n2039), .B2(n2061), .ZN(n3400)
         );
  OAI22_X1 U1272 ( .A1(n6559), .A2(n6653), .B1(n2039), .B2(n2060), .ZN(n3401)
         );
  OAI22_X1 U1273 ( .A1(n6585), .A2(n6641), .B1(n6584), .B2(n2031), .ZN(n3493)
         );
  OAI22_X1 U1274 ( .A1(n6586), .A2(n6644), .B1(n2010), .B2(n2030), .ZN(n3494)
         );
  OAI22_X1 U1275 ( .A1(n6586), .A2(n6647), .B1(n6584), .B2(n2029), .ZN(n3495)
         );
  OAI22_X1 U1276 ( .A1(n6586), .A2(n6650), .B1(n2010), .B2(n2028), .ZN(n3496)
         );
  OAI22_X1 U1277 ( .A1(n6586), .A2(n6656), .B1(n6584), .B2(n2027), .ZN(n3498)
         );
  OAI22_X1 U1278 ( .A1(n6587), .A2(n6659), .B1(n2010), .B2(n2026), .ZN(n3499)
         );
  OAI22_X1 U1279 ( .A1(n6587), .A2(n6662), .B1(n2010), .B2(n2025), .ZN(n3500)
         );
  OAI22_X1 U1280 ( .A1(n6594), .A2(n6635), .B1(n6593), .B2(n2006), .ZN(n3523)
         );
  OAI22_X1 U1281 ( .A1(n6594), .A2(n6638), .B1(n1978), .B2(n2005), .ZN(n3524)
         );
  OAI22_X1 U1282 ( .A1(n6594), .A2(n6641), .B1(n6593), .B2(n2004), .ZN(n3525)
         );
  OAI22_X1 U1283 ( .A1(n6595), .A2(n6644), .B1(n1978), .B2(n2003), .ZN(n3526)
         );
  OAI22_X1 U1284 ( .A1(n6595), .A2(n6647), .B1(n6593), .B2(n2002), .ZN(n3527)
         );
  OAI22_X1 U1285 ( .A1(n6595), .A2(n6650), .B1(n1978), .B2(n2001), .ZN(n3528)
         );
  OAI22_X1 U1286 ( .A1(n6595), .A2(n6653), .B1(n1978), .B2(n2000), .ZN(n3529)
         );
  OAI22_X1 U1287 ( .A1(n6621), .A2(n6641), .B1(n6620), .B2(n1964), .ZN(n3621)
         );
  OAI22_X1 U1288 ( .A1(n6622), .A2(n6644), .B1(n6620), .B2(n1963), .ZN(n3622)
         );
  OAI22_X1 U1289 ( .A1(n6622), .A2(n6647), .B1(n6620), .B2(n1962), .ZN(n3623)
         );
  OAI22_X1 U1290 ( .A1(n6622), .A2(n6650), .B1(n6620), .B2(n1961), .ZN(n3624)
         );
  OAI22_X1 U1291 ( .A1(n6622), .A2(n6656), .B1(n6620), .B2(n1960), .ZN(n3626)
         );
  OAI22_X1 U1292 ( .A1(n6623), .A2(n6659), .B1(n1944), .B2(n1959), .ZN(n3627)
         );
  OAI22_X1 U1293 ( .A1(n6623), .A2(n6662), .B1(n1944), .B2(n1958), .ZN(n3628)
         );
  OAI22_X1 U1294 ( .A1(n6723), .A2(n6635), .B1(n6722), .B2(n1937), .ZN(n3651)
         );
  OAI22_X1 U1295 ( .A1(n6723), .A2(n6638), .B1(n1880), .B2(n1935), .ZN(n3652)
         );
  OAI22_X1 U1296 ( .A1(n6723), .A2(n6641), .B1(n6722), .B2(n1933), .ZN(n3653)
         );
  OAI22_X1 U1297 ( .A1(n6724), .A2(n6644), .B1(n1880), .B2(n1931), .ZN(n3654)
         );
  OAI22_X1 U1298 ( .A1(n6724), .A2(n6647), .B1(n6722), .B2(n1929), .ZN(n3655)
         );
  OAI22_X1 U1299 ( .A1(n6724), .A2(n6650), .B1(n1880), .B2(n1927), .ZN(n3656)
         );
  OAI22_X1 U1300 ( .A1(n6724), .A2(n6653), .B1(n1880), .B2(n1925), .ZN(n3657)
         );
  OAI22_X1 U1301 ( .A1(n6405), .A2(n6629), .B1(n6404), .B2(n2332), .ZN(n2849)
         );
  OAI22_X1 U1302 ( .A1(n6407), .A2(n6670), .B1(n6404), .B2(n2323), .ZN(n2862)
         );
  OAI22_X1 U1303 ( .A1(n6407), .A2(n6673), .B1(n6404), .B2(n2322), .ZN(n2863)
         );
  OAI22_X1 U1304 ( .A1(n6408), .A2(n6676), .B1(n6404), .B2(n2321), .ZN(n2864)
         );
  OAI22_X1 U1305 ( .A1(n6408), .A2(n6679), .B1(n6404), .B2(n2320), .ZN(n2865)
         );
  OAI22_X1 U1306 ( .A1(n6408), .A2(n6682), .B1(n6404), .B2(n2319), .ZN(n2866)
         );
  OAI22_X1 U1307 ( .A1(n6408), .A2(n6685), .B1(n6404), .B2(n2318), .ZN(n2867)
         );
  OAI22_X1 U1308 ( .A1(n6408), .A2(n6688), .B1(n6404), .B2(n2317), .ZN(n2868)
         );
  OAI22_X1 U1309 ( .A1(n6409), .A2(n6691), .B1(n6404), .B2(n2316), .ZN(n2869)
         );
  OAI22_X1 U1310 ( .A1(n6409), .A2(n6694), .B1(n6404), .B2(n2315), .ZN(n2870)
         );
  OAI22_X1 U1311 ( .A1(n6409), .A2(n6697), .B1(n6404), .B2(n2314), .ZN(n2871)
         );
  OAI22_X1 U1312 ( .A1(n6409), .A2(n6700), .B1(n6404), .B2(n2313), .ZN(n2872)
         );
  OAI22_X1 U1313 ( .A1(n6409), .A2(n6703), .B1(n6404), .B2(n2312), .ZN(n2873)
         );
  OAI22_X1 U1314 ( .A1(n6415), .A2(n6658), .B1(n6413), .B2(n2299), .ZN(n2890)
         );
  OAI22_X1 U1315 ( .A1(n6416), .A2(n6670), .B1(n6413), .B2(n2298), .ZN(n2894)
         );
  OAI22_X1 U1316 ( .A1(n6416), .A2(n6673), .B1(n6413), .B2(n2297), .ZN(n2895)
         );
  OAI22_X1 U1317 ( .A1(n6417), .A2(n6676), .B1(n6413), .B2(n2296), .ZN(n2896)
         );
  OAI22_X1 U1318 ( .A1(n6417), .A2(n6679), .B1(n6413), .B2(n2295), .ZN(n2897)
         );
  OAI22_X1 U1319 ( .A1(n6417), .A2(n6682), .B1(n6413), .B2(n2294), .ZN(n2898)
         );
  OAI22_X1 U1320 ( .A1(n6417), .A2(n6685), .B1(n6413), .B2(n2293), .ZN(n2899)
         );
  OAI22_X1 U1321 ( .A1(n6417), .A2(n6688), .B1(n6413), .B2(n2292), .ZN(n2900)
         );
  OAI22_X1 U1322 ( .A1(n6418), .A2(n6691), .B1(n6413), .B2(n2291), .ZN(n2901)
         );
  OAI22_X1 U1323 ( .A1(n6418), .A2(n6694), .B1(n6413), .B2(n2290), .ZN(n2902)
         );
  OAI22_X1 U1324 ( .A1(n6418), .A2(n6697), .B1(n6413), .B2(n2289), .ZN(n2903)
         );
  OAI22_X1 U1325 ( .A1(n6418), .A2(n6703), .B1(n6413), .B2(n2287), .ZN(n2905)
         );
  OAI22_X1 U1326 ( .A1(n6420), .A2(n6733), .B1(n6413), .B2(n2280), .ZN(n2912)
         );
  OAI22_X1 U1327 ( .A1(n6442), .A2(n6657), .B1(n6440), .B2(n2265), .ZN(n2986)
         );
  OAI22_X1 U1328 ( .A1(n6443), .A2(n6669), .B1(n6440), .B2(n2264), .ZN(n2990)
         );
  OAI22_X1 U1329 ( .A1(n6443), .A2(n6672), .B1(n6440), .B2(n2263), .ZN(n2991)
         );
  OAI22_X1 U1330 ( .A1(n6444), .A2(n6675), .B1(n6440), .B2(n2262), .ZN(n2992)
         );
  OAI22_X1 U1331 ( .A1(n6444), .A2(n6678), .B1(n6440), .B2(n2261), .ZN(n2993)
         );
  OAI22_X1 U1332 ( .A1(n6444), .A2(n6681), .B1(n6440), .B2(n2260), .ZN(n2994)
         );
  OAI22_X1 U1333 ( .A1(n6444), .A2(n6684), .B1(n6440), .B2(n2259), .ZN(n2995)
         );
  OAI22_X1 U1334 ( .A1(n6444), .A2(n6687), .B1(n6440), .B2(n2258), .ZN(n2996)
         );
  OAI22_X1 U1335 ( .A1(n6445), .A2(n6690), .B1(n6440), .B2(n2257), .ZN(n2997)
         );
  OAI22_X1 U1336 ( .A1(n6445), .A2(n6693), .B1(n6440), .B2(n2256), .ZN(n2998)
         );
  OAI22_X1 U1337 ( .A1(n6445), .A2(n6696), .B1(n6440), .B2(n2255), .ZN(n2999)
         );
  OAI22_X1 U1338 ( .A1(n6445), .A2(n6702), .B1(n6440), .B2(n2253), .ZN(n3001)
         );
  OAI22_X1 U1339 ( .A1(n6447), .A2(n6732), .B1(n6440), .B2(n2246), .ZN(n3008)
         );
  OAI22_X1 U1340 ( .A1(n6450), .A2(n6629), .B1(n6449), .B2(n2242), .ZN(n3009)
         );
  OAI22_X1 U1341 ( .A1(n6452), .A2(n6669), .B1(n6449), .B2(n2233), .ZN(n3022)
         );
  OAI22_X1 U1342 ( .A1(n6452), .A2(n6672), .B1(n6449), .B2(n2232), .ZN(n3023)
         );
  OAI22_X1 U1343 ( .A1(n6453), .A2(n6675), .B1(n6449), .B2(n2231), .ZN(n3024)
         );
  OAI22_X1 U1344 ( .A1(n6453), .A2(n6678), .B1(n6449), .B2(n2230), .ZN(n3025)
         );
  OAI22_X1 U1345 ( .A1(n6453), .A2(n6681), .B1(n6449), .B2(n2229), .ZN(n3026)
         );
  OAI22_X1 U1346 ( .A1(n6453), .A2(n6684), .B1(n6449), .B2(n2228), .ZN(n3027)
         );
  OAI22_X1 U1347 ( .A1(n6453), .A2(n6687), .B1(n6449), .B2(n2227), .ZN(n3028)
         );
  OAI22_X1 U1348 ( .A1(n6454), .A2(n6690), .B1(n6449), .B2(n2226), .ZN(n3029)
         );
  OAI22_X1 U1349 ( .A1(n6454), .A2(n6693), .B1(n6449), .B2(n2225), .ZN(n3030)
         );
  OAI22_X1 U1350 ( .A1(n6454), .A2(n6696), .B1(n6449), .B2(n2224), .ZN(n3031)
         );
  OAI22_X1 U1351 ( .A1(n6454), .A2(n6699), .B1(n6449), .B2(n2223), .ZN(n3032)
         );
  OAI22_X1 U1352 ( .A1(n6454), .A2(n6702), .B1(n6449), .B2(n2222), .ZN(n3033)
         );
  OAI22_X1 U1353 ( .A1(n6478), .A2(n6657), .B1(n6476), .B2(n2205), .ZN(n3114)
         );
  OAI22_X1 U1354 ( .A1(n6479), .A2(n6669), .B1(n6476), .B2(n2204), .ZN(n3118)
         );
  OAI22_X1 U1355 ( .A1(n6479), .A2(n6672), .B1(n6476), .B2(n2203), .ZN(n3119)
         );
  OAI22_X1 U1356 ( .A1(n6480), .A2(n6675), .B1(n6476), .B2(n2202), .ZN(n3120)
         );
  OAI22_X1 U1357 ( .A1(n6480), .A2(n6678), .B1(n6476), .B2(n2201), .ZN(n3121)
         );
  OAI22_X1 U1358 ( .A1(n6480), .A2(n6681), .B1(n6476), .B2(n2200), .ZN(n3122)
         );
  OAI22_X1 U1359 ( .A1(n6480), .A2(n6684), .B1(n6476), .B2(n2199), .ZN(n3123)
         );
  OAI22_X1 U1360 ( .A1(n6480), .A2(n6687), .B1(n6476), .B2(n2198), .ZN(n3124)
         );
  OAI22_X1 U1361 ( .A1(n6481), .A2(n6690), .B1(n6476), .B2(n2197), .ZN(n3125)
         );
  OAI22_X1 U1362 ( .A1(n6481), .A2(n6693), .B1(n6476), .B2(n2196), .ZN(n3126)
         );
  OAI22_X1 U1363 ( .A1(n6481), .A2(n6696), .B1(n6476), .B2(n2195), .ZN(n3127)
         );
  OAI22_X1 U1364 ( .A1(n6481), .A2(n6702), .B1(n6476), .B2(n2193), .ZN(n3129)
         );
  OAI22_X1 U1365 ( .A1(n6483), .A2(n6732), .B1(n6476), .B2(n2186), .ZN(n3136)
         );
  OAI22_X1 U1366 ( .A1(n6486), .A2(n6630), .B1(n6485), .B2(n2182), .ZN(n3137)
         );
  OAI22_X1 U1367 ( .A1(n6488), .A2(n6669), .B1(n6485), .B2(n2173), .ZN(n3150)
         );
  OAI22_X1 U1368 ( .A1(n6488), .A2(n6672), .B1(n6485), .B2(n2172), .ZN(n3151)
         );
  OAI22_X1 U1369 ( .A1(n6489), .A2(n6675), .B1(n6485), .B2(n2171), .ZN(n3152)
         );
  OAI22_X1 U1370 ( .A1(n6489), .A2(n6678), .B1(n6485), .B2(n2170), .ZN(n3153)
         );
  OAI22_X1 U1371 ( .A1(n6489), .A2(n6681), .B1(n6485), .B2(n2169), .ZN(n3154)
         );
  OAI22_X1 U1372 ( .A1(n6489), .A2(n6684), .B1(n6485), .B2(n2168), .ZN(n3155)
         );
  OAI22_X1 U1373 ( .A1(n6489), .A2(n6687), .B1(n6485), .B2(n2167), .ZN(n3156)
         );
  OAI22_X1 U1374 ( .A1(n6490), .A2(n6690), .B1(n6485), .B2(n2166), .ZN(n3157)
         );
  OAI22_X1 U1375 ( .A1(n6490), .A2(n6693), .B1(n6485), .B2(n2165), .ZN(n3158)
         );
  OAI22_X1 U1376 ( .A1(n6490), .A2(n6696), .B1(n6485), .B2(n2164), .ZN(n3159)
         );
  OAI22_X1 U1377 ( .A1(n6490), .A2(n6699), .B1(n6485), .B2(n2163), .ZN(n3160)
         );
  OAI22_X1 U1378 ( .A1(n6490), .A2(n6702), .B1(n6485), .B2(n2162), .ZN(n3161)
         );
  OAI22_X1 U1379 ( .A1(n6513), .A2(n6630), .B1(n6512), .B2(n2153), .ZN(n3233)
         );
  OAI22_X1 U1380 ( .A1(n6515), .A2(n6669), .B1(n6512), .B2(n2144), .ZN(n3246)
         );
  OAI22_X1 U1381 ( .A1(n6515), .A2(n6672), .B1(n6512), .B2(n2143), .ZN(n3247)
         );
  OAI22_X1 U1382 ( .A1(n6516), .A2(n6675), .B1(n6512), .B2(n2142), .ZN(n3248)
         );
  OAI22_X1 U1383 ( .A1(n6516), .A2(n6678), .B1(n6512), .B2(n2141), .ZN(n3249)
         );
  OAI22_X1 U1384 ( .A1(n6516), .A2(n6681), .B1(n6512), .B2(n2140), .ZN(n3250)
         );
  OAI22_X1 U1385 ( .A1(n6516), .A2(n6684), .B1(n6512), .B2(n2139), .ZN(n3251)
         );
  OAI22_X1 U1386 ( .A1(n6516), .A2(n6687), .B1(n6512), .B2(n2138), .ZN(n3252)
         );
  OAI22_X1 U1387 ( .A1(n6517), .A2(n6690), .B1(n6512), .B2(n2137), .ZN(n3253)
         );
  OAI22_X1 U1388 ( .A1(n6517), .A2(n6693), .B1(n6512), .B2(n2136), .ZN(n3254)
         );
  OAI22_X1 U1389 ( .A1(n6517), .A2(n6696), .B1(n6512), .B2(n2135), .ZN(n3255)
         );
  OAI22_X1 U1390 ( .A1(n6517), .A2(n6699), .B1(n6512), .B2(n2134), .ZN(n3256)
         );
  OAI22_X1 U1391 ( .A1(n6517), .A2(n6702), .B1(n6512), .B2(n2133), .ZN(n3257)
         );
  OAI22_X1 U1392 ( .A1(n6523), .A2(n6657), .B1(n6521), .B2(n2120), .ZN(n3274)
         );
  OAI22_X1 U1393 ( .A1(n6524), .A2(n6669), .B1(n6521), .B2(n2119), .ZN(n3278)
         );
  OAI22_X1 U1394 ( .A1(n6524), .A2(n6672), .B1(n6521), .B2(n2118), .ZN(n3279)
         );
  OAI22_X1 U1395 ( .A1(n6525), .A2(n6675), .B1(n6521), .B2(n2117), .ZN(n3280)
         );
  OAI22_X1 U1396 ( .A1(n6525), .A2(n6678), .B1(n6521), .B2(n2116), .ZN(n3281)
         );
  OAI22_X1 U1397 ( .A1(n6525), .A2(n6681), .B1(n6521), .B2(n2115), .ZN(n3282)
         );
  OAI22_X1 U1398 ( .A1(n6525), .A2(n6684), .B1(n6521), .B2(n2114), .ZN(n3283)
         );
  OAI22_X1 U1399 ( .A1(n6525), .A2(n6687), .B1(n6521), .B2(n2113), .ZN(n3284)
         );
  OAI22_X1 U1400 ( .A1(n6526), .A2(n6690), .B1(n6521), .B2(n2112), .ZN(n3285)
         );
  OAI22_X1 U1401 ( .A1(n6526), .A2(n6693), .B1(n6521), .B2(n2111), .ZN(n3286)
         );
  OAI22_X1 U1402 ( .A1(n6526), .A2(n6696), .B1(n6521), .B2(n2110), .ZN(n3287)
         );
  OAI22_X1 U1403 ( .A1(n6526), .A2(n6702), .B1(n6521), .B2(n2108), .ZN(n3289)
         );
  OAI22_X1 U1404 ( .A1(n6528), .A2(n6732), .B1(n6521), .B2(n2101), .ZN(n3296)
         );
  OAI22_X1 U1405 ( .A1(n6549), .A2(n6630), .B1(n6548), .B2(n2094), .ZN(n3361)
         );
  OAI22_X1 U1406 ( .A1(n6551), .A2(n6662), .B1(n6548), .B2(n2085), .ZN(n3372)
         );
  OAI22_X1 U1407 ( .A1(n6551), .A2(n6665), .B1(n6548), .B2(n2084), .ZN(n3373)
         );
  OAI22_X1 U1408 ( .A1(n6551), .A2(n6668), .B1(n6548), .B2(n2083), .ZN(n3374)
         );
  OAI22_X1 U1409 ( .A1(n6551), .A2(n6671), .B1(n6548), .B2(n2082), .ZN(n3375)
         );
  OAI22_X1 U1410 ( .A1(n6552), .A2(n6674), .B1(n6548), .B2(n2081), .ZN(n3376)
         );
  OAI22_X1 U1411 ( .A1(n6552), .A2(n6677), .B1(n6548), .B2(n2080), .ZN(n3377)
         );
  OAI22_X1 U1412 ( .A1(n6552), .A2(n6680), .B1(n6548), .B2(n2079), .ZN(n3378)
         );
  OAI22_X1 U1413 ( .A1(n6552), .A2(n6683), .B1(n6548), .B2(n2078), .ZN(n3379)
         );
  OAI22_X1 U1414 ( .A1(n6552), .A2(n6686), .B1(n6548), .B2(n2077), .ZN(n3380)
         );
  OAI22_X1 U1415 ( .A1(n6553), .A2(n6689), .B1(n6548), .B2(n2076), .ZN(n3381)
         );
  OAI22_X1 U1416 ( .A1(n6553), .A2(n6692), .B1(n6548), .B2(n2075), .ZN(n3382)
         );
  OAI22_X1 U1417 ( .A1(n6553), .A2(n6695), .B1(n6548), .B2(n2074), .ZN(n3383)
         );
  OAI22_X1 U1418 ( .A1(n6559), .A2(n6656), .B1(n6557), .B2(n2059), .ZN(n3402)
         );
  OAI22_X1 U1419 ( .A1(n6560), .A2(n6668), .B1(n6557), .B2(n2058), .ZN(n3406)
         );
  OAI22_X1 U1420 ( .A1(n6560), .A2(n6671), .B1(n6557), .B2(n2057), .ZN(n3407)
         );
  OAI22_X1 U1421 ( .A1(n6561), .A2(n6674), .B1(n6557), .B2(n2056), .ZN(n3408)
         );
  OAI22_X1 U1422 ( .A1(n6561), .A2(n6677), .B1(n6557), .B2(n2055), .ZN(n3409)
         );
  OAI22_X1 U1423 ( .A1(n6561), .A2(n6680), .B1(n6557), .B2(n2054), .ZN(n3410)
         );
  OAI22_X1 U1424 ( .A1(n6561), .A2(n6683), .B1(n6557), .B2(n2053), .ZN(n3411)
         );
  OAI22_X1 U1425 ( .A1(n6561), .A2(n6686), .B1(n6557), .B2(n2052), .ZN(n3412)
         );
  OAI22_X1 U1426 ( .A1(n6562), .A2(n6689), .B1(n6557), .B2(n2051), .ZN(n3413)
         );
  OAI22_X1 U1427 ( .A1(n6562), .A2(n6692), .B1(n6557), .B2(n2050), .ZN(n3414)
         );
  OAI22_X1 U1428 ( .A1(n6562), .A2(n6695), .B1(n6557), .B2(n2049), .ZN(n3415)
         );
  OAI22_X1 U1429 ( .A1(n6562), .A2(n6701), .B1(n6557), .B2(n2047), .ZN(n3417)
         );
  OAI22_X1 U1430 ( .A1(n6564), .A2(n6731), .B1(n6557), .B2(n2040), .ZN(n3424)
         );
  OAI22_X1 U1431 ( .A1(n6585), .A2(n6631), .B1(n6584), .B2(n2033), .ZN(n3489)
         );
  OAI22_X1 U1432 ( .A1(n6587), .A2(n6665), .B1(n6584), .B2(n2024), .ZN(n3501)
         );
  OAI22_X1 U1433 ( .A1(n6587), .A2(n6668), .B1(n6584), .B2(n2023), .ZN(n3502)
         );
  OAI22_X1 U1434 ( .A1(n6587), .A2(n6671), .B1(n6584), .B2(n2022), .ZN(n3503)
         );
  OAI22_X1 U1435 ( .A1(n6588), .A2(n6674), .B1(n6584), .B2(n2021), .ZN(n3504)
         );
  OAI22_X1 U1436 ( .A1(n6588), .A2(n6677), .B1(n6584), .B2(n2020), .ZN(n3505)
         );
  OAI22_X1 U1437 ( .A1(n6588), .A2(n6680), .B1(n6584), .B2(n2019), .ZN(n3506)
         );
  OAI22_X1 U1438 ( .A1(n6588), .A2(n6683), .B1(n6584), .B2(n2018), .ZN(n3507)
         );
  OAI22_X1 U1439 ( .A1(n6588), .A2(n6686), .B1(n6584), .B2(n2017), .ZN(n3508)
         );
  OAI22_X1 U1440 ( .A1(n6589), .A2(n6689), .B1(n6584), .B2(n2016), .ZN(n3509)
         );
  OAI22_X1 U1441 ( .A1(n6589), .A2(n6692), .B1(n6584), .B2(n2015), .ZN(n3510)
         );
  OAI22_X1 U1442 ( .A1(n6589), .A2(n6695), .B1(n6584), .B2(n2014), .ZN(n3511)
         );
  OAI22_X1 U1443 ( .A1(n6589), .A2(n6698), .B1(n6584), .B2(n2013), .ZN(n3512)
         );
  OAI22_X1 U1444 ( .A1(n6595), .A2(n6656), .B1(n6593), .B2(n1999), .ZN(n3530)
         );
  OAI22_X1 U1445 ( .A1(n6596), .A2(n6665), .B1(n6593), .B2(n1998), .ZN(n3533)
         );
  OAI22_X1 U1446 ( .A1(n6596), .A2(n6668), .B1(n6593), .B2(n1997), .ZN(n3534)
         );
  OAI22_X1 U1447 ( .A1(n6596), .A2(n6671), .B1(n6593), .B2(n1996), .ZN(n3535)
         );
  OAI22_X1 U1448 ( .A1(n6597), .A2(n6674), .B1(n6593), .B2(n1995), .ZN(n3536)
         );
  OAI22_X1 U1449 ( .A1(n6597), .A2(n6677), .B1(n6593), .B2(n1994), .ZN(n3537)
         );
  OAI22_X1 U1450 ( .A1(n6597), .A2(n6680), .B1(n6593), .B2(n1993), .ZN(n3538)
         );
  OAI22_X1 U1451 ( .A1(n6597), .A2(n6683), .B1(n6593), .B2(n1992), .ZN(n3539)
         );
  OAI22_X1 U1452 ( .A1(n6597), .A2(n6686), .B1(n6593), .B2(n1991), .ZN(n3540)
         );
  OAI22_X1 U1453 ( .A1(n6598), .A2(n6689), .B1(n6593), .B2(n1990), .ZN(n3541)
         );
  OAI22_X1 U1454 ( .A1(n6598), .A2(n6692), .B1(n6593), .B2(n1989), .ZN(n3542)
         );
  OAI22_X1 U1455 ( .A1(n6598), .A2(n6695), .B1(n6593), .B2(n1988), .ZN(n3543)
         );
  OAI22_X1 U1456 ( .A1(n6600), .A2(n6731), .B1(n6593), .B2(n1979), .ZN(n3552)
         );
  OAI22_X1 U1457 ( .A1(n6621), .A2(n6631), .B1(n6620), .B2(n1966), .ZN(n3617)
         );
  OAI22_X1 U1458 ( .A1(n6623), .A2(n6665), .B1(n6620), .B2(n1957), .ZN(n3629)
         );
  OAI22_X1 U1459 ( .A1(n6623), .A2(n6668), .B1(n6620), .B2(n1956), .ZN(n3630)
         );
  OAI22_X1 U1460 ( .A1(n6623), .A2(n6671), .B1(n6620), .B2(n1955), .ZN(n3631)
         );
  OAI22_X1 U1461 ( .A1(n6624), .A2(n6674), .B1(n6620), .B2(n1954), .ZN(n3632)
         );
  OAI22_X1 U1462 ( .A1(n6624), .A2(n6677), .B1(n6620), .B2(n1953), .ZN(n3633)
         );
  OAI22_X1 U1463 ( .A1(n6624), .A2(n6680), .B1(n6620), .B2(n1952), .ZN(n3634)
         );
  OAI22_X1 U1464 ( .A1(n6624), .A2(n6683), .B1(n6620), .B2(n1951), .ZN(n3635)
         );
  OAI22_X1 U1465 ( .A1(n6624), .A2(n6686), .B1(n6620), .B2(n1950), .ZN(n3636)
         );
  OAI22_X1 U1466 ( .A1(n6625), .A2(n6689), .B1(n6620), .B2(n1949), .ZN(n3637)
         );
  OAI22_X1 U1467 ( .A1(n6625), .A2(n6692), .B1(n6620), .B2(n1948), .ZN(n3638)
         );
  OAI22_X1 U1468 ( .A1(n6625), .A2(n6695), .B1(n6620), .B2(n1947), .ZN(n3639)
         );
  OAI22_X1 U1469 ( .A1(n6625), .A2(n6698), .B1(n6620), .B2(n1946), .ZN(n3640)
         );
  OAI22_X1 U1470 ( .A1(n6724), .A2(n6656), .B1(n6722), .B2(n1923), .ZN(n3658)
         );
  OAI22_X1 U1471 ( .A1(n6725), .A2(n6665), .B1(n6722), .B2(n1919), .ZN(n3661)
         );
  OAI22_X1 U1472 ( .A1(n6725), .A2(n6668), .B1(n6722), .B2(n1917), .ZN(n3662)
         );
  OAI22_X1 U1473 ( .A1(n6725), .A2(n6671), .B1(n6722), .B2(n1915), .ZN(n3663)
         );
  OAI22_X1 U1474 ( .A1(n6726), .A2(n6674), .B1(n6722), .B2(n1913), .ZN(n3664)
         );
  OAI22_X1 U1475 ( .A1(n6726), .A2(n6677), .B1(n6722), .B2(n1911), .ZN(n3665)
         );
  OAI22_X1 U1476 ( .A1(n6726), .A2(n6680), .B1(n6722), .B2(n1909), .ZN(n3666)
         );
  OAI22_X1 U1477 ( .A1(n6726), .A2(n6683), .B1(n6722), .B2(n1907), .ZN(n3667)
         );
  OAI22_X1 U1478 ( .A1(n6726), .A2(n6686), .B1(n6722), .B2(n1905), .ZN(n3668)
         );
  OAI22_X1 U1479 ( .A1(n6727), .A2(n6689), .B1(n6722), .B2(n1903), .ZN(n3669)
         );
  OAI22_X1 U1480 ( .A1(n6727), .A2(n6692), .B1(n6722), .B2(n1901), .ZN(n3670)
         );
  OAI22_X1 U1481 ( .A1(n6727), .A2(n6695), .B1(n6722), .B2(n1899), .ZN(n3671)
         );
  OAI22_X1 U1482 ( .A1(n6729), .A2(n6731), .B1(n6722), .B2(n1881), .ZN(n3680)
         );
  OAI22_X1 U1483 ( .A1(n6405), .A2(n6634), .B1(n2310), .B2(n2331), .ZN(n2850)
         );
  OAI22_X1 U1484 ( .A1(n6410), .A2(n6706), .B1(n6404), .B2(n2311), .ZN(n2874)
         );
  OAI22_X1 U1485 ( .A1(n6450), .A2(n6633), .B1(n2220), .B2(n2241), .ZN(n3010)
         );
  OAI22_X1 U1486 ( .A1(n6455), .A2(n6705), .B1(n6449), .B2(n2221), .ZN(n3034)
         );
  OAI22_X1 U1487 ( .A1(n6486), .A2(n6633), .B1(n2160), .B2(n2181), .ZN(n3138)
         );
  OAI22_X1 U1488 ( .A1(n6491), .A2(n6705), .B1(n6485), .B2(n2161), .ZN(n3162)
         );
  OAI22_X1 U1489 ( .A1(n6513), .A2(n6633), .B1(n2131), .B2(n2152), .ZN(n3234)
         );
  OAI22_X1 U1490 ( .A1(n6518), .A2(n6705), .B1(n6512), .B2(n2132), .ZN(n3258)
         );
  OAI22_X1 U1491 ( .A1(n6621), .A2(n6632), .B1(n1944), .B2(n1965), .ZN(n3618)
         );
  OAI22_X1 U1492 ( .A1(n6625), .A2(n6701), .B1(n6620), .B2(n1945), .ZN(n3641)
         );
  OAI22_X1 U1493 ( .A1(n6585), .A2(n6632), .B1(n2010), .B2(n2032), .ZN(n3490)
         );
  OAI22_X1 U1494 ( .A1(n6589), .A2(n6701), .B1(n2010), .B2(n2012), .ZN(n3513)
         );
  OAI22_X1 U1495 ( .A1(n6590), .A2(n6704), .B1(n6584), .B2(n2011), .ZN(n3514)
         );
  OAI22_X1 U1496 ( .A1(n6549), .A2(n6632), .B1(n2070), .B2(n2093), .ZN(n3362)
         );
  OAI22_X1 U1497 ( .A1(n6553), .A2(n6698), .B1(n2070), .B2(n2073), .ZN(n3384)
         );
  OAI22_X1 U1498 ( .A1(n6553), .A2(n6701), .B1(n2070), .B2(n2072), .ZN(n3385)
         );
  OAI22_X1 U1499 ( .A1(n6554), .A2(n6704), .B1(n6548), .B2(n2071), .ZN(n3386)
         );
  OAI22_X1 U1500 ( .A1(n6414), .A2(n6634), .B1(n2279), .B2(n2307), .ZN(n2882)
         );
  OAI22_X1 U1501 ( .A1(n6418), .A2(n6700), .B1(n2279), .B2(n2288), .ZN(n2904)
         );
  OAI22_X1 U1502 ( .A1(n6419), .A2(n6706), .B1(n2279), .B2(n2286), .ZN(n2906)
         );
  OAI22_X1 U1503 ( .A1(n6419), .A2(n6709), .B1(n2279), .B2(n2285), .ZN(n2907)
         );
  OAI22_X1 U1504 ( .A1(n6419), .A2(n6712), .B1(n2279), .B2(n2284), .ZN(n2908)
         );
  OAI22_X1 U1505 ( .A1(n6419), .A2(n6715), .B1(n2279), .B2(n2283), .ZN(n2909)
         );
  OAI22_X1 U1506 ( .A1(n6419), .A2(n6718), .B1(n2279), .B2(n2282), .ZN(n2910)
         );
  OAI22_X1 U1507 ( .A1(n6420), .A2(n6721), .B1(n6413), .B2(n2281), .ZN(n2911)
         );
  OAI22_X1 U1508 ( .A1(n6441), .A2(n6633), .B1(n2245), .B2(n2273), .ZN(n2978)
         );
  OAI22_X1 U1509 ( .A1(n6445), .A2(n6699), .B1(n2245), .B2(n2254), .ZN(n3000)
         );
  OAI22_X1 U1510 ( .A1(n6446), .A2(n6705), .B1(n2245), .B2(n2252), .ZN(n3002)
         );
  OAI22_X1 U1511 ( .A1(n6446), .A2(n6708), .B1(n2245), .B2(n2251), .ZN(n3003)
         );
  OAI22_X1 U1512 ( .A1(n6446), .A2(n6711), .B1(n2245), .B2(n2250), .ZN(n3004)
         );
  OAI22_X1 U1513 ( .A1(n6446), .A2(n6714), .B1(n2245), .B2(n2249), .ZN(n3005)
         );
  OAI22_X1 U1514 ( .A1(n6446), .A2(n6717), .B1(n2245), .B2(n2248), .ZN(n3006)
         );
  OAI22_X1 U1515 ( .A1(n6447), .A2(n6720), .B1(n6440), .B2(n2247), .ZN(n3007)
         );
  OAI22_X1 U1516 ( .A1(n6477), .A2(n6633), .B1(n2185), .B2(n2213), .ZN(n3106)
         );
  OAI22_X1 U1517 ( .A1(n6481), .A2(n6699), .B1(n2185), .B2(n2194), .ZN(n3128)
         );
  OAI22_X1 U1518 ( .A1(n6482), .A2(n6705), .B1(n2185), .B2(n2192), .ZN(n3130)
         );
  OAI22_X1 U1519 ( .A1(n6482), .A2(n6708), .B1(n2185), .B2(n2191), .ZN(n3131)
         );
  OAI22_X1 U1520 ( .A1(n6482), .A2(n6711), .B1(n2185), .B2(n2190), .ZN(n3132)
         );
  OAI22_X1 U1521 ( .A1(n6482), .A2(n6714), .B1(n2185), .B2(n2189), .ZN(n3133)
         );
  OAI22_X1 U1522 ( .A1(n6482), .A2(n6717), .B1(n2185), .B2(n2188), .ZN(n3134)
         );
  OAI22_X1 U1523 ( .A1(n6483), .A2(n6720), .B1(n6476), .B2(n2187), .ZN(n3135)
         );
  OAI22_X1 U1524 ( .A1(n6522), .A2(n6633), .B1(n2100), .B2(n2128), .ZN(n3266)
         );
  OAI22_X1 U1525 ( .A1(n6526), .A2(n6699), .B1(n2100), .B2(n2109), .ZN(n3288)
         );
  OAI22_X1 U1526 ( .A1(n6527), .A2(n6705), .B1(n2100), .B2(n2107), .ZN(n3290)
         );
  OAI22_X1 U1527 ( .A1(n6527), .A2(n6708), .B1(n2100), .B2(n2106), .ZN(n3291)
         );
  OAI22_X1 U1528 ( .A1(n6527), .A2(n6711), .B1(n2100), .B2(n2105), .ZN(n3292)
         );
  OAI22_X1 U1529 ( .A1(n6527), .A2(n6714), .B1(n2100), .B2(n2104), .ZN(n3293)
         );
  OAI22_X1 U1530 ( .A1(n6527), .A2(n6717), .B1(n2100), .B2(n2103), .ZN(n3294)
         );
  OAI22_X1 U1531 ( .A1(n6528), .A2(n6720), .B1(n6521), .B2(n2102), .ZN(n3295)
         );
  OAI22_X1 U1532 ( .A1(n6558), .A2(n6632), .B1(n2039), .B2(n2067), .ZN(n3394)
         );
  OAI22_X1 U1533 ( .A1(n6562), .A2(n6698), .B1(n2039), .B2(n2048), .ZN(n3416)
         );
  OAI22_X1 U1534 ( .A1(n6563), .A2(n6704), .B1(n2039), .B2(n2046), .ZN(n3418)
         );
  OAI22_X1 U1535 ( .A1(n6563), .A2(n6707), .B1(n2039), .B2(n2045), .ZN(n3419)
         );
  OAI22_X1 U1536 ( .A1(n6563), .A2(n6710), .B1(n2039), .B2(n2044), .ZN(n3420)
         );
  OAI22_X1 U1537 ( .A1(n6563), .A2(n6713), .B1(n2039), .B2(n2043), .ZN(n3421)
         );
  OAI22_X1 U1538 ( .A1(n6563), .A2(n6716), .B1(n2039), .B2(n2042), .ZN(n3422)
         );
  OAI22_X1 U1539 ( .A1(n6564), .A2(n6719), .B1(n6557), .B2(n2041), .ZN(n3423)
         );
  OAI22_X1 U1540 ( .A1(n6594), .A2(n6632), .B1(n1978), .B2(n2007), .ZN(n3522)
         );
  OAI22_X1 U1541 ( .A1(n6598), .A2(n6698), .B1(n1978), .B2(n1987), .ZN(n3544)
         );
  OAI22_X1 U1542 ( .A1(n6598), .A2(n6701), .B1(n1978), .B2(n1986), .ZN(n3545)
         );
  OAI22_X1 U1543 ( .A1(n6599), .A2(n6704), .B1(n1978), .B2(n1985), .ZN(n3546)
         );
  OAI22_X1 U1544 ( .A1(n6599), .A2(n6707), .B1(n1978), .B2(n1984), .ZN(n3547)
         );
  OAI22_X1 U1545 ( .A1(n6599), .A2(n6710), .B1(n1978), .B2(n1983), .ZN(n3548)
         );
  OAI22_X1 U1546 ( .A1(n6599), .A2(n6713), .B1(n6593), .B2(n1982), .ZN(n3549)
         );
  OAI22_X1 U1547 ( .A1(n6599), .A2(n6716), .B1(n1978), .B2(n1981), .ZN(n3550)
         );
  OAI22_X1 U1548 ( .A1(n6600), .A2(n6719), .B1(n6593), .B2(n1980), .ZN(n3551)
         );
  OAI22_X1 U1549 ( .A1(n6723), .A2(n6632), .B1(n1880), .B2(n1939), .ZN(n3650)
         );
  OAI22_X1 U1550 ( .A1(n6727), .A2(n6698), .B1(n1880), .B2(n1897), .ZN(n3672)
         );
  OAI22_X1 U1551 ( .A1(n6727), .A2(n6701), .B1(n1880), .B2(n1895), .ZN(n3673)
         );
  OAI22_X1 U1552 ( .A1(n6728), .A2(n6704), .B1(n1880), .B2(n1893), .ZN(n3674)
         );
  OAI22_X1 U1553 ( .A1(n6728), .A2(n6707), .B1(n1880), .B2(n1891), .ZN(n3675)
         );
  OAI22_X1 U1554 ( .A1(n6728), .A2(n6710), .B1(n1880), .B2(n1889), .ZN(n3676)
         );
  OAI22_X1 U1555 ( .A1(n6728), .A2(n6713), .B1(n6722), .B2(n1887), .ZN(n3677)
         );
  OAI22_X1 U1556 ( .A1(n6728), .A2(n6716), .B1(n1880), .B2(n1885), .ZN(n3678)
         );
  OAI22_X1 U1557 ( .A1(n6729), .A2(n6719), .B1(n6722), .B2(n1883), .ZN(n3679)
         );
  NAND2_X1 U1558 ( .A1(DATAIN[20]), .A2(n6734), .ZN(n1902) );
  NAND2_X1 U1559 ( .A1(DATAIN[21]), .A2(n6734), .ZN(n1900) );
  NAND2_X1 U1560 ( .A1(DATAIN[22]), .A2(n6734), .ZN(n1898) );
  NAND2_X1 U1561 ( .A1(DATAIN[23]), .A2(n6734), .ZN(n1896) );
  NAND2_X1 U1562 ( .A1(DATAIN[24]), .A2(n6734), .ZN(n1894) );
  NAND2_X1 U1563 ( .A1(DATAIN[25]), .A2(n6734), .ZN(n1892) );
  NAND2_X1 U1564 ( .A1(DATAIN[26]), .A2(n6734), .ZN(n1890) );
  NAND2_X1 U1565 ( .A1(DATAIN[27]), .A2(n6734), .ZN(n1888) );
  NAND2_X1 U1566 ( .A1(DATAIN[28]), .A2(n6734), .ZN(n1886) );
  NAND2_X1 U1567 ( .A1(DATAIN[29]), .A2(n6734), .ZN(n1884) );
  NAND2_X1 U1568 ( .A1(DATAIN[30]), .A2(n6734), .ZN(n1882) );
  NAND2_X1 U1569 ( .A1(DATAIN[31]), .A2(n6734), .ZN(n1879) );
  AND2_X1 U1570 ( .A1(n5051), .A2(n5059), .ZN(n2378) );
  AND2_X1 U1571 ( .A1(n5045), .A2(n5058), .ZN(n2373) );
  AND2_X1 U1572 ( .A1(n5045), .A2(n5059), .ZN(n2371) );
  AND2_X1 U1573 ( .A1(n5058), .A2(n5051), .ZN(n2380) );
  AND2_X1 U1574 ( .A1(n5070), .A2(n5051), .ZN(n2398) );
  AND2_X1 U1575 ( .A1(n5071), .A2(n5051), .ZN(n2396) );
  AND2_X1 U1576 ( .A1(n5079), .A2(n5051), .ZN(n2405) );
  AND2_X1 U1577 ( .A1(n5080), .A2(n5051), .ZN(n2403) );
  AND2_X1 U1578 ( .A1(n5070), .A2(n5045), .ZN(n2391) );
  AND2_X1 U1579 ( .A1(n5071), .A2(n5045), .ZN(n2389) );
  AND2_X1 U1580 ( .A1(n5079), .A2(n5045), .ZN(n2410) );
  NAND2_X1 U1581 ( .A1(DATAIN[8]), .A2(n6734), .ZN(n1924) );
  NAND2_X1 U1582 ( .A1(DATAIN[9]), .A2(n6735), .ZN(n1922) );
  NAND2_X1 U1583 ( .A1(DATAIN[10]), .A2(n6734), .ZN(n1921) );
  NAND2_X1 U1584 ( .A1(DATAIN[11]), .A2(n6735), .ZN(n1920) );
  NAND2_X1 U1585 ( .A1(DATAIN[12]), .A2(n6734), .ZN(n1918) );
  NAND2_X1 U1586 ( .A1(DATAIN[13]), .A2(n6734), .ZN(n1916) );
  NAND2_X1 U1587 ( .A1(DATAIN[14]), .A2(n6734), .ZN(n1914) );
  NAND2_X1 U1588 ( .A1(DATAIN[15]), .A2(n6734), .ZN(n1912) );
  NAND2_X1 U1589 ( .A1(DATAIN[16]), .A2(n6734), .ZN(n1910) );
  NAND2_X1 U1590 ( .A1(DATAIN[17]), .A2(n6734), .ZN(n1908) );
  NAND2_X1 U1591 ( .A1(DATAIN[18]), .A2(n6734), .ZN(n1906) );
  NAND2_X1 U1592 ( .A1(DATAIN[19]), .A2(n6735), .ZN(n1904) );
  NAND2_X1 U1593 ( .A1(DATAIN[0]), .A2(n6735), .ZN(n1940) );
  NAND2_X1 U1594 ( .A1(DATAIN[1]), .A2(n6735), .ZN(n1938) );
  NAND2_X1 U1595 ( .A1(DATAIN[2]), .A2(n6734), .ZN(n1936) );
  NAND2_X1 U1596 ( .A1(DATAIN[3]), .A2(n6734), .ZN(n1934) );
  NAND2_X1 U1597 ( .A1(DATAIN[4]), .A2(n6734), .ZN(n1932) );
  NAND2_X1 U1598 ( .A1(DATAIN[5]), .A2(n6735), .ZN(n1930) );
  NAND2_X1 U1599 ( .A1(DATAIN[6]), .A2(n6734), .ZN(n1928) );
  NAND2_X1 U1600 ( .A1(DATAIN[7]), .A2(n6735), .ZN(n1926) );
  OAI21_X1 U1601 ( .B1(n1973), .B2(n2339), .A(n6735), .ZN(n2346) );
  INV_X1 U1602 ( .A(n1972), .ZN(n6610) );
  OAI21_X1 U1603 ( .B1(n1941), .B2(n1973), .A(RESET), .ZN(n1972) );
  INV_X1 U1604 ( .A(n2336), .ZN(n6394) );
  OAI21_X1 U1605 ( .B1(n1973), .B2(n2308), .A(RESET), .ZN(n2336) );
  INV_X1 U1606 ( .A(n2277), .ZN(n6430) );
  OAI21_X1 U1607 ( .B1(n1973), .B2(n2243), .A(RESET), .ZN(n2277) );
  INV_X1 U1608 ( .A(n2217), .ZN(n6466) );
  OAI21_X1 U1609 ( .B1(n1973), .B2(n2183), .A(RESET), .ZN(n2217) );
  INV_X1 U1610 ( .A(n2157), .ZN(n6502) );
  OAI21_X1 U1611 ( .B1(n1973), .B2(n2129), .A(RESET), .ZN(n2157) );
  INV_X1 U1612 ( .A(n2098), .ZN(n6538) );
  OAI21_X1 U1613 ( .B1(n1973), .B2(n2068), .A(n6735), .ZN(n2098) );
  INV_X1 U1614 ( .A(n2037), .ZN(n6574) );
  OAI21_X1 U1615 ( .B1(n1973), .B2(n2008), .A(n6735), .ZN(n2037) );
  INV_X1 U1616 ( .A(n2343), .ZN(n6376) );
  OAI21_X1 U1617 ( .B1(n1967), .B2(n2339), .A(n6735), .ZN(n2343) );
  INV_X1 U1618 ( .A(n2310), .ZN(n6412) );
  OAI21_X1 U1619 ( .B1(n1967), .B2(n2308), .A(RESET), .ZN(n2310) );
  INV_X1 U1620 ( .A(n2245), .ZN(n6448) );
  OAI21_X1 U1621 ( .B1(n1967), .B2(n2243), .A(RESET), .ZN(n2245) );
  INV_X1 U1622 ( .A(n2185), .ZN(n6484) );
  OAI21_X1 U1623 ( .B1(n1967), .B2(n2183), .A(RESET), .ZN(n2185) );
  INV_X1 U1624 ( .A(n2131), .ZN(n6520) );
  OAI21_X1 U1625 ( .B1(n1967), .B2(n2129), .A(RESET), .ZN(n2131) );
  INV_X1 U1626 ( .A(n2070), .ZN(n6556) );
  OAI21_X1 U1627 ( .B1(n1967), .B2(n2068), .A(RESET), .ZN(n2070) );
  INV_X1 U1628 ( .A(n2010), .ZN(n6592) );
  OAI21_X1 U1629 ( .B1(n1967), .B2(n2008), .A(RESET), .ZN(n2010) );
  INV_X1 U1630 ( .A(n2334), .ZN(n6403) );
  OAI21_X1 U1631 ( .B1(n1970), .B2(n2308), .A(RESET), .ZN(n2334) );
  INV_X1 U1632 ( .A(n2279), .ZN(n6421) );
  OAI21_X1 U1633 ( .B1(n1942), .B2(n2308), .A(RESET), .ZN(n2279) );
  INV_X1 U1634 ( .A(n2275), .ZN(n6439) );
  OAI21_X1 U1635 ( .B1(n1970), .B2(n2243), .A(RESET), .ZN(n2275) );
  INV_X1 U1636 ( .A(n2220), .ZN(n6457) );
  OAI21_X1 U1637 ( .B1(n1942), .B2(n2243), .A(RESET), .ZN(n2220) );
  INV_X1 U1638 ( .A(n2215), .ZN(n6475) );
  OAI21_X1 U1639 ( .B1(n1970), .B2(n2183), .A(RESET), .ZN(n2215) );
  NOR3_X1 U1640 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n5695) );
  NOR3_X1 U1641 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n5691), .ZN(n5694) );
  NOR3_X1 U1642 ( .A1(n5691), .A2(ADD_RD1[3]), .A3(n5705), .ZN(n5703) );
  NOR3_X1 U1643 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n5705), .ZN(n5702) );
  NOR3_X1 U1644 ( .A1(n5692), .A2(ADD_RD1[0]), .A3(n5705), .ZN(n5707) );
  OAI221_X1 U1645 ( .B1(n448), .B2(n5982), .C1(n2242), .C2(n5991), .A(n5701), 
        .ZN(n5700) );
  AOI22_X1 U1646 ( .A1(n5997), .A2(n5068), .B1(n6005), .B2(n5069), .ZN(n5701)
         );
  OAI221_X1 U1647 ( .B1(n445), .B2(n6097), .C1(n2153), .C2(n6106), .A(n5683), 
        .ZN(n5682) );
  AOI22_X1 U1648 ( .A1(n6112), .A2(n5042), .B1(n6114), .B2(n5043), .ZN(n5683)
         );
  OAI221_X1 U1649 ( .B1(n441), .B2(n5982), .C1(n2236), .C2(n5990), .A(n5673), 
        .ZN(n5672) );
  AOI22_X1 U1650 ( .A1(n5997), .A2(n5024), .B1(n6005), .B2(n5025), .ZN(n5673)
         );
  OAI221_X1 U1651 ( .B1(n438), .B2(n6097), .C1(n2147), .C2(n6106), .A(n5665), 
        .ZN(n5664) );
  AOI22_X1 U1652 ( .A1(n6113), .A2(n5008), .B1(n6115), .B2(n5009), .ZN(n5665)
         );
  OAI221_X1 U1653 ( .B1(n434), .B2(n5983), .C1(n2235), .C2(n5990), .A(n5655), 
        .ZN(n5654) );
  AOI22_X1 U1654 ( .A1(n5997), .A2(n4990), .B1(n6005), .B2(n4991), .ZN(n5655)
         );
  OAI221_X1 U1655 ( .B1(n431), .B2(n6100), .C1(n2146), .C2(n6107), .A(n5647), 
        .ZN(n5646) );
  AOI22_X1 U1656 ( .A1(n5096), .A2(n4974), .B1(n5097), .B2(n4975), .ZN(n5647)
         );
  OAI221_X1 U1657 ( .B1(n427), .B2(n5983), .C1(n2234), .C2(n5992), .A(n5637), 
        .ZN(n5636) );
  AOI22_X1 U1658 ( .A1(n5998), .A2(n4956), .B1(n6006), .B2(n4957), .ZN(n5637)
         );
  OAI221_X1 U1659 ( .B1(n424), .B2(n6098), .C1(n2145), .C2(n6107), .A(n5629), 
        .ZN(n5628) );
  AOI22_X1 U1660 ( .A1(n6112), .A2(n4940), .B1(n6114), .B2(n4941), .ZN(n5629)
         );
  OAI221_X1 U1661 ( .B1(n2265), .B2(n5983), .C1(n7), .C2(n5991), .A(n5119), 
        .ZN(n5116) );
  AOI22_X1 U1662 ( .A1(n6000), .A2(n2390), .B1(n6010), .B2(n2392), .ZN(n5119)
         );
  OAI221_X1 U1663 ( .B1(n2120), .B2(n6098), .C1(n4), .C2(n6109), .A(n5095), 
        .ZN(n5092) );
  AOI22_X1 U1664 ( .A1(n6113), .A2(n2358), .B1(n6115), .B2(n2360), .ZN(n5095)
         );
  OAI221_X1 U1665 ( .B1(n2246), .B2(n5986), .C1(n56), .C2(n5995), .A(n5259), 
        .ZN(n5258) );
  AOI22_X1 U1666 ( .A1(n5997), .A2(n2641), .B1(n6005), .B2(n2642), .ZN(n5259)
         );
  OAI221_X1 U1667 ( .B1(n2101), .B2(n6102), .C1(n53), .C2(n6110), .A(n5251), 
        .ZN(n5250) );
  AOI22_X1 U1668 ( .A1(n6112), .A2(n2625), .B1(n6114), .B2(n2626), .ZN(n5251)
         );
  OAI221_X1 U1669 ( .B1(n2271), .B2(n5984), .C1(n49), .C2(n5991), .A(n5241), 
        .ZN(n5240) );
  AOI22_X1 U1670 ( .A1(n5998), .A2(n2607), .B1(n6006), .B2(n2608), .ZN(n5241)
         );
  OAI221_X1 U1671 ( .B1(n2126), .B2(n6102), .C1(n46), .C2(n6110), .A(n5233), 
        .ZN(n5232) );
  AOI22_X1 U1672 ( .A1(n6113), .A2(n2591), .B1(n6115), .B2(n2592), .ZN(n5233)
         );
  OAI221_X1 U1673 ( .B1(n2270), .B2(n5987), .C1(n42), .C2(n5995), .A(n5223), 
        .ZN(n5222) );
  AOI22_X1 U1674 ( .A1(n6002), .A2(n2573), .B1(n6007), .B2(n2574), .ZN(n5223)
         );
  OAI221_X1 U1675 ( .B1(n2125), .B2(n6103), .C1(n39), .C2(n6111), .A(n5215), 
        .ZN(n5214) );
  AOI22_X1 U1676 ( .A1(n5096), .A2(n2557), .B1(n5097), .B2(n2558), .ZN(n5215)
         );
  OAI221_X1 U1677 ( .B1(n2251), .B2(n5986), .C1(n98), .C2(n5990), .A(n5367), 
        .ZN(n5366) );
  AOI22_X1 U1678 ( .A1(n6003), .A2(n4446), .B1(n6011), .B2(n4447), .ZN(n5367)
         );
  OAI221_X1 U1679 ( .B1(n2106), .B2(n6098), .C1(n95), .C2(n6110), .A(n5359), 
        .ZN(n5358) );
  AOI22_X1 U1680 ( .A1(n6112), .A2(n4430), .B1(n6114), .B2(n4431), .ZN(n5359)
         );
  OAI221_X1 U1681 ( .B1(n2250), .B2(n5987), .C1(n91), .C2(n5994), .A(n5349), 
        .ZN(n5348) );
  AOI22_X1 U1682 ( .A1(n6002), .A2(n4412), .B1(n6011), .B2(n4413), .ZN(n5349)
         );
  OAI221_X1 U1683 ( .B1(n2105), .B2(n6101), .C1(n88), .C2(n6109), .A(n5341), 
        .ZN(n5340) );
  AOI22_X1 U1684 ( .A1(n6113), .A2(n4396), .B1(n6115), .B2(n4397), .ZN(n5341)
         );
  OAI221_X1 U1685 ( .B1(n2249), .B2(n5986), .C1(n84), .C2(n5994), .A(n5331), 
        .ZN(n5330) );
  AOI22_X1 U1686 ( .A1(n6001), .A2(n4378), .B1(n6006), .B2(n4379), .ZN(n5331)
         );
  OAI221_X1 U1687 ( .B1(n2104), .B2(n6102), .C1(n81), .C2(n6110), .A(n5323), 
        .ZN(n5322) );
  AOI22_X1 U1688 ( .A1(n5096), .A2(n4362), .B1(n5097), .B2(n4363), .ZN(n5323)
         );
  OAI221_X1 U1689 ( .B1(n2248), .B2(n5986), .C1(n77), .C2(n5994), .A(n5313), 
        .ZN(n5312) );
  AOI22_X1 U1690 ( .A1(n6000), .A2(n4344), .B1(n6007), .B2(n4345), .ZN(n5313)
         );
  OAI221_X1 U1691 ( .B1(n2103), .B2(n6103), .C1(n74), .C2(n6110), .A(n5305), 
        .ZN(n5304) );
  AOI22_X1 U1692 ( .A1(n6112), .A2(n4328), .B1(n6114), .B2(n4329), .ZN(n5305)
         );
  OAI221_X1 U1693 ( .B1(n2272), .B2(n5987), .C1(n70), .C2(n5995), .A(n5295), 
        .ZN(n5294) );
  AOI22_X1 U1694 ( .A1(n5997), .A2(n4310), .B1(n6005), .B2(n4311), .ZN(n5295)
         );
  OAI221_X1 U1695 ( .B1(n2127), .B2(n6102), .C1(n67), .C2(n6111), .A(n5287), 
        .ZN(n5286) );
  AOI22_X1 U1696 ( .A1(n6113), .A2(n3718), .B1(n6115), .B2(n3719), .ZN(n5287)
         );
  OAI221_X1 U1697 ( .B1(n2247), .B2(n5987), .C1(n63), .C2(n5995), .A(n5277), 
        .ZN(n5276) );
  AOI22_X1 U1698 ( .A1(n6002), .A2(n3700), .B1(n6011), .B2(n3701), .ZN(n5277)
         );
  OAI221_X1 U1699 ( .B1(n2102), .B2(n6103), .C1(n60), .C2(n6111), .A(n5269), 
        .ZN(n5268) );
  AOI22_X1 U1700 ( .A1(n5096), .A2(n3684), .B1(n5097), .B2(n3685), .ZN(n5269)
         );
  OAI221_X1 U1701 ( .B1(n447), .B2(n5950), .C1(n2182), .C2(n5959), .A(n5704), 
        .ZN(n5699) );
  AOI22_X1 U1702 ( .A1(n5965), .A2(n5073), .B1(n5973), .B2(n5074), .ZN(n5704)
         );
  OAI221_X1 U1703 ( .B1(n440), .B2(n5950), .C1(n2176), .C2(n5958), .A(n5674), 
        .ZN(n5671) );
  AOI22_X1 U1704 ( .A1(n5965), .A2(n5027), .B1(n5973), .B2(n5028), .ZN(n5674)
         );
  OAI221_X1 U1705 ( .B1(n433), .B2(n5951), .C1(n2175), .C2(n5958), .A(n5656), 
        .ZN(n5653) );
  AOI22_X1 U1706 ( .A1(n5965), .A2(n4993), .B1(n5973), .B2(n4994), .ZN(n5656)
         );
  OAI221_X1 U1707 ( .B1(n426), .B2(n5951), .C1(n2174), .C2(n5960), .A(n5638), 
        .ZN(n5635) );
  AOI22_X1 U1708 ( .A1(n5966), .A2(n4959), .B1(n5974), .B2(n4960), .ZN(n5638)
         );
  OAI221_X1 U1709 ( .B1(n423), .B2(n6082), .C1(n2084), .C2(n6087), .A(n5630), 
        .ZN(n5627) );
  AOI22_X1 U1710 ( .A1(n6092), .A2(n4943), .B1(n6094), .B2(n4944), .ZN(n5630)
         );
  OAI221_X1 U1711 ( .B1(n2205), .B2(n5951), .C1(n6), .C2(n5959), .A(n5124), 
        .ZN(n5115) );
  AOI22_X1 U1712 ( .A1(n5968), .A2(n2397), .B1(n5978), .B2(n2399), .ZN(n5124)
         );
  OAI221_X1 U1713 ( .B1(n2186), .B2(n5954), .C1(n55), .C2(n5963), .A(n5260), 
        .ZN(n5257) );
  AOI22_X1 U1714 ( .A1(n5965), .A2(n2644), .B1(n5973), .B2(n2645), .ZN(n5260)
         );
  OAI221_X1 U1715 ( .B1(n2211), .B2(n5952), .C1(n48), .C2(n5959), .A(n5242), 
        .ZN(n5239) );
  AOI22_X1 U1716 ( .A1(n5966), .A2(n2610), .B1(n5974), .B2(n2611), .ZN(n5242)
         );
  OAI221_X1 U1717 ( .B1(n2210), .B2(n5955), .C1(n41), .C2(n5963), .A(n5224), 
        .ZN(n5221) );
  AOI22_X1 U1718 ( .A1(n5970), .A2(n2576), .B1(n5975), .B2(n2577), .ZN(n5224)
         );
  OAI221_X1 U1719 ( .B1(n2191), .B2(n5954), .C1(n97), .C2(n5958), .A(n5368), 
        .ZN(n5365) );
  AOI22_X1 U1720 ( .A1(n5971), .A2(n4449), .B1(n5979), .B2(n4450), .ZN(n5368)
         );
  OAI221_X1 U1721 ( .B1(n2045), .B2(n6082), .C1(n94), .C2(n6090), .A(n5360), 
        .ZN(n5357) );
  AOI22_X1 U1722 ( .A1(n6092), .A2(n4433), .B1(n6094), .B2(n4434), .ZN(n5360)
         );
  OAI221_X1 U1723 ( .B1(n2190), .B2(n5955), .C1(n90), .C2(n5962), .A(n5350), 
        .ZN(n5347) );
  AOI22_X1 U1724 ( .A1(n5970), .A2(n4415), .B1(n5979), .B2(n4416), .ZN(n5350)
         );
  OAI221_X1 U1725 ( .B1(n2044), .B2(n6078), .C1(n87), .C2(n6091), .A(n5342), 
        .ZN(n5339) );
  AOI22_X1 U1726 ( .A1(n6093), .A2(n4399), .B1(n6095), .B2(n4400), .ZN(n5342)
         );
  OAI221_X1 U1727 ( .B1(n2189), .B2(n5954), .C1(n83), .C2(n5962), .A(n5332), 
        .ZN(n5329) );
  AOI22_X1 U1728 ( .A1(n5969), .A2(n4381), .B1(n5974), .B2(n4382), .ZN(n5332)
         );
  OAI221_X1 U1729 ( .B1(n2043), .B2(n6082), .C1(n80), .C2(n6090), .A(n5324), 
        .ZN(n5321) );
  AOI22_X1 U1730 ( .A1(n5101), .A2(n4365), .B1(n5102), .B2(n4366), .ZN(n5324)
         );
  OAI221_X1 U1731 ( .B1(n2188), .B2(n5954), .C1(n76), .C2(n5962), .A(n5314), 
        .ZN(n5311) );
  AOI22_X1 U1732 ( .A1(n5968), .A2(n4347), .B1(n5975), .B2(n4348), .ZN(n5314)
         );
  OAI221_X1 U1733 ( .B1(n2042), .B2(n6083), .C1(n73), .C2(n6090), .A(n5306), 
        .ZN(n5303) );
  AOI22_X1 U1734 ( .A1(n6092), .A2(n4331), .B1(n6094), .B2(n4332), .ZN(n5306)
         );
  OAI221_X1 U1735 ( .B1(n2212), .B2(n5955), .C1(n69), .C2(n5963), .A(n5296), 
        .ZN(n5293) );
  AOI22_X1 U1736 ( .A1(n5965), .A2(n4313), .B1(n5973), .B2(n4314), .ZN(n5296)
         );
  OAI221_X1 U1737 ( .B1(n2187), .B2(n5955), .C1(n62), .C2(n5963), .A(n5278), 
        .ZN(n5275) );
  AOI22_X1 U1738 ( .A1(n5970), .A2(n3703), .B1(n5979), .B2(n3704), .ZN(n5278)
         );
  OAI221_X1 U1739 ( .B1(n446), .B2(n5922), .C1(n2332), .C2(n5925), .A(n5706), 
        .ZN(n5698) );
  AOI22_X1 U1740 ( .A1(n5933), .A2(n5077), .B1(n5941), .B2(n5078), .ZN(n5706)
         );
  OAI221_X1 U1741 ( .B1(n443), .B2(n6045), .C1(n2033), .C2(n6053), .A(n5693), 
        .ZN(n5680) );
  AOI22_X1 U1742 ( .A1(n6061), .A2(n5056), .B1(n6070), .B2(n5057), .ZN(n5693)
         );
  OAI221_X1 U1743 ( .B1(n439), .B2(n5918), .C1(n2326), .C2(n5926), .A(n5675), 
        .ZN(n5670) );
  AOI22_X1 U1744 ( .A1(n5933), .A2(n5030), .B1(n5941), .B2(n5031), .ZN(n5675)
         );
  OAI221_X1 U1745 ( .B1(n436), .B2(n6045), .C1(n2026), .C2(n6057), .A(n5667), 
        .ZN(n5662) );
  AOI22_X1 U1746 ( .A1(n6061), .A2(n5014), .B1(n6070), .B2(n5015), .ZN(n5667)
         );
  OAI221_X1 U1747 ( .B1(n432), .B2(n5919), .C1(n2325), .C2(n5926), .A(n5657), 
        .ZN(n5652) );
  AOI22_X1 U1748 ( .A1(n5933), .A2(n4996), .B1(n5941), .B2(n4997), .ZN(n5657)
         );
  OAI221_X1 U1749 ( .B1(n429), .B2(n6050), .C1(n2025), .C2(n6059), .A(n5649), 
        .ZN(n5644) );
  AOI22_X1 U1750 ( .A1(n6061), .A2(n4980), .B1(n6070), .B2(n4981), .ZN(n5649)
         );
  OAI221_X1 U1751 ( .B1(n425), .B2(n5919), .C1(n2324), .C2(n5929), .A(n5639), 
        .ZN(n5634) );
  AOI22_X1 U1752 ( .A1(n5934), .A2(n4962), .B1(n5942), .B2(n4963), .ZN(n5639)
         );
  OAI221_X1 U1753 ( .B1(n4079), .B2(n5891), .C1(n4078), .C2(n5895), .A(n5478), 
        .ZN(n5471) );
  AOI22_X1 U1754 ( .A1(n5907), .A2(n4659), .B1(n5915), .B2(n4660), .ZN(n5478)
         );
  OAI221_X1 U1755 ( .B1(n4061), .B2(n5888), .C1(n4060), .C2(n5897), .A(n5460), 
        .ZN(n5453) );
  AOI22_X1 U1756 ( .A1(n5907), .A2(n4625), .B1(n5915), .B2(n4626), .ZN(n5460)
         );
  OAI221_X1 U1757 ( .B1(n4043), .B2(n5886), .C1(n4042), .C2(n5896), .A(n5442), 
        .ZN(n5435) );
  AOI22_X1 U1758 ( .A1(n5906), .A2(n4591), .B1(n5912), .B2(n4592), .ZN(n5442)
         );
  OAI221_X1 U1759 ( .B1(n4025), .B2(n5887), .C1(n4024), .C2(n5897), .A(n5424), 
        .ZN(n5417) );
  AOI22_X1 U1760 ( .A1(n5906), .A2(n4557), .B1(n5914), .B2(n4558), .ZN(n5424)
         );
  OAI221_X1 U1761 ( .B1(n4151), .B2(n5887), .C1(n4150), .C2(n5896), .A(n5550), 
        .ZN(n5543) );
  AOI22_X1 U1762 ( .A1(n5904), .A2(n4795), .B1(n5912), .B2(n4796), .ZN(n5550)
         );
  OAI221_X1 U1763 ( .B1(n4133), .B2(n5889), .C1(n4132), .C2(n5896), .A(n5532), 
        .ZN(n5525) );
  AOI22_X1 U1764 ( .A1(n5903), .A2(n4761), .B1(n5913), .B2(n4762), .ZN(n5532)
         );
  OAI221_X1 U1765 ( .B1(n4115), .B2(n5888), .C1(n4114), .C2(n5898), .A(n5514), 
        .ZN(n5507) );
  AOI22_X1 U1766 ( .A1(n5906), .A2(n4727), .B1(n5914), .B2(n4728), .ZN(n5514)
         );
  OAI221_X1 U1767 ( .B1(n4097), .B2(n5889), .C1(n4096), .C2(n5894), .A(n5496), 
        .ZN(n5489) );
  AOI22_X1 U1768 ( .A1(n5906), .A2(n4693), .B1(n5914), .B2(n4694), .ZN(n5496)
         );
  OAI221_X1 U1769 ( .B1(n4223), .B2(n5885), .C1(n4222), .C2(n5895), .A(n5622), 
        .ZN(n5615) );
  AOI22_X1 U1771 ( .A1(n5904), .A2(n4931), .B1(n5911), .B2(n4932), .ZN(n5622)
         );
  OAI221_X1 U1772 ( .B1(n4205), .B2(n5887), .C1(n4204), .C2(n5895), .A(n5604), 
        .ZN(n5597) );
  AOI22_X1 U1774 ( .A1(n5903), .A2(n4897), .B1(n5911), .B2(n4898), .ZN(n5604)
         );
  OAI221_X1 U1775 ( .B1(n4187), .B2(n5890), .C1(n4186), .C2(n5896), .A(n5586), 
        .ZN(n5579) );
  AOI22_X1 U1776 ( .A1(n5902), .A2(n4863), .B1(n5912), .B2(n4864), .ZN(n5586)
         );
  OAI221_X1 U1777 ( .B1(n4169), .B2(n5887), .C1(n4168), .C2(n5897), .A(n5568), 
        .ZN(n5561) );
  AOI22_X1 U1779 ( .A1(n5905), .A2(n4829), .B1(n5913), .B2(n4830), .ZN(n5568)
         );
  OAI221_X1 U1780 ( .B1(n4295), .B2(n5885), .C1(n4294), .C2(n5895), .A(n5711), 
        .ZN(n5697) );
  AOI22_X1 U1781 ( .A1(n5902), .A2(n5084), .B1(n5910), .B2(n5085), .ZN(n5711)
         );
  OAI221_X1 U1782 ( .B1(n442), .B2(n6018), .C1(n1966), .C2(n6021), .A(n5696), 
        .ZN(n5679) );
  AOI22_X1 U1784 ( .A1(n6030), .A2(n5061), .B1(n6037), .B2(n5062), .ZN(n5696)
         );
  OAI221_X1 U1785 ( .B1(n4277), .B2(n5885), .C1(n4276), .C2(n5897), .A(n5676), 
        .ZN(n5669) );
  AOI22_X1 U1786 ( .A1(n5902), .A2(n5033), .B1(n5910), .B2(n5034), .ZN(n5676)
         );
  OAI221_X1 U1787 ( .B1(n435), .B2(n6014), .C1(n1959), .C2(n6021), .A(n5668), 
        .ZN(n5661) );
  AOI22_X1 U1788 ( .A1(n6030), .A2(n5017), .B1(n6037), .B2(n5018), .ZN(n5668)
         );
  OAI221_X1 U1789 ( .B1(n4259), .B2(n5886), .C1(n4258), .C2(n5894), .A(n5658), 
        .ZN(n5651) );
  AOI22_X1 U1790 ( .A1(n5903), .A2(n4999), .B1(n5910), .B2(n5000), .ZN(n5658)
         );
  OAI221_X1 U1791 ( .B1(n428), .B2(n6019), .C1(n1958), .C2(n6022), .A(n5650), 
        .ZN(n5643) );
  AOI22_X1 U1792 ( .A1(n6030), .A2(n4983), .B1(n6037), .B2(n4984), .ZN(n5650)
         );
  OAI221_X1 U1793 ( .B1(n4241), .B2(n5886), .C1(n4240), .C2(n5894), .A(n5640), 
        .ZN(n5633) );
  AOI22_X1 U1794 ( .A1(n5903), .A2(n4965), .B1(n5911), .B2(n4966), .ZN(n5640)
         );
  OAI221_X1 U1795 ( .B1(n3791), .B2(n5885), .C1(n3790), .C2(n5896), .A(n5190), 
        .ZN(n5183) );
  AOI22_X1 U1796 ( .A1(n5905), .A2(n2514), .B1(n5912), .B2(n2515), .ZN(n5190)
         );
  OAI221_X1 U1797 ( .B1(n3773), .B2(n5886), .C1(n3772), .C2(n5895), .A(n5172), 
        .ZN(n5165) );
  AOI22_X1 U1798 ( .A1(n5905), .A2(n2480), .B1(n5913), .B2(n2481), .ZN(n5172)
         );
  OAI221_X1 U1799 ( .B1(n3755), .B2(n5886), .C1(n3754), .C2(n5894), .A(n5154), 
        .ZN(n5147) );
  AOI22_X1 U1800 ( .A1(n5905), .A2(n2446), .B1(n5913), .B2(n2447), .ZN(n5154)
         );
  OAI221_X1 U1801 ( .B1(n3737), .B2(n5890), .C1(n3736), .C2(n5894), .A(n5134), 
        .ZN(n5113) );
  AOI22_X1 U1802 ( .A1(n5906), .A2(n2411), .B1(n5914), .B2(n2413), .ZN(n5134)
         );
  OAI221_X1 U1803 ( .B1(n3863), .B2(n5891), .C1(n3862), .C2(n5899), .A(n5262), 
        .ZN(n5255) );
  AOI22_X1 U1804 ( .A1(n5905), .A2(n2650), .B1(n5910), .B2(n2651), .ZN(n5262)
         );
  OAI221_X1 U1805 ( .B1(n3845), .B2(n5891), .C1(n3844), .C2(n5898), .A(n5244), 
        .ZN(n5237) );
  AOI22_X1 U1806 ( .A1(n5903), .A2(n2616), .B1(n5911), .B2(n2617), .ZN(n5244)
         );
  OAI221_X1 U1807 ( .B1(n3827), .B2(n5890), .C1(n3826), .C2(n5899), .A(n5226), 
        .ZN(n5219) );
  AOI22_X1 U1808 ( .A1(n5904), .A2(n2582), .B1(n5911), .B2(n2583), .ZN(n5226)
         );
  OAI221_X1 U1809 ( .B1(n3809), .B2(n5889), .C1(n3808), .C2(n5899), .A(n5208), 
        .ZN(n5201) );
  AOI22_X1 U1810 ( .A1(n5904), .A2(n2548), .B1(n5914), .B2(n2549), .ZN(n5208)
         );
  OAI221_X1 U1811 ( .B1(n4007), .B2(n5887), .C1(n4006), .C2(n5897), .A(n5406), 
        .ZN(n5399) );
  AOI22_X1 U1812 ( .A1(n5907), .A2(n4523), .B1(n5915), .B2(n4524), .ZN(n5406)
         );
  OAI221_X1 U1813 ( .B1(n3989), .B2(n5890), .C1(n3988), .C2(n5897), .A(n5388), 
        .ZN(n5381) );
  AOI22_X1 U1814 ( .A1(n5907), .A2(n4489), .B1(n5913), .B2(n4490), .ZN(n5388)
         );
  OAI221_X1 U1815 ( .B1(n3971), .B2(n5888), .C1(n3970), .C2(n5898), .A(n5370), 
        .ZN(n5363) );
  AOI22_X1 U1816 ( .A1(n5906), .A2(n4455), .B1(n5915), .B2(n4456), .ZN(n5370)
         );
  OAI221_X1 U1817 ( .B1(n3953), .B2(n5889), .C1(n3952), .C2(n5894), .A(n5352), 
        .ZN(n5345) );
  AOI22_X1 U1818 ( .A1(n5906), .A2(n4421), .B1(n5914), .B2(n4422), .ZN(n5352)
         );
  OAI221_X1 U1819 ( .B1(n3935), .B2(n5888), .C1(n3934), .C2(n5898), .A(n5334), 
        .ZN(n5327) );
  AOI22_X1 U1820 ( .A1(n5902), .A2(n4387), .B1(n5915), .B2(n4388), .ZN(n5334)
         );
  OAI221_X1 U1821 ( .B1(n3917), .B2(n5891), .C1(n3916), .C2(n5898), .A(n5316), 
        .ZN(n5309) );
  AOI22_X1 U1822 ( .A1(n5902), .A2(n4353), .B1(n5915), .B2(n4354), .ZN(n5316)
         );
  OAI221_X1 U1823 ( .B1(n3899), .B2(n5890), .C1(n3898), .C2(n5899), .A(n5298), 
        .ZN(n5291) );
  AOI22_X1 U1824 ( .A1(n5902), .A2(n4319), .B1(n5910), .B2(n4320), .ZN(n5298)
         );
  OAI221_X1 U1825 ( .B1(n3881), .B2(n5890), .C1(n3880), .C2(n5899), .A(n5280), 
        .ZN(n5273) );
  AOI22_X1 U1826 ( .A1(n5907), .A2(n3709), .B1(n5914), .B2(n3710), .ZN(n5280)
         );
  OAI221_X1 U1827 ( .B1(n2000), .B2(n6046), .C1(n9), .C2(n6054), .A(n5145), 
        .ZN(n5140) );
  AOI22_X1 U1828 ( .A1(n6063), .A2(n2427), .B1(n6073), .B2(n2428), .ZN(n5145)
         );
  OAI221_X1 U1829 ( .B1(n2299), .B2(n5918), .C1(n5), .C2(n5929), .A(n5129), 
        .ZN(n5114) );
  AOI22_X1 U1830 ( .A1(n5936), .A2(n2404), .B1(n5946), .B2(n2406), .ZN(n5129)
         );
  OAI221_X1 U1831 ( .B1(n2280), .B2(n5923), .C1(n54), .C2(n5931), .A(n5261), 
        .ZN(n5256) );
  AOI22_X1 U1832 ( .A1(n5933), .A2(n2647), .B1(n5941), .B2(n2648), .ZN(n5261)
         );
  OAI221_X1 U1833 ( .B1(n1979), .B2(n6051), .C1(n51), .C2(n6058), .A(n5253), 
        .ZN(n5248) );
  AOI22_X1 U1834 ( .A1(n6061), .A2(n2631), .B1(n6070), .B2(n2632), .ZN(n5253)
         );
  OAI221_X1 U1835 ( .B1(n2305), .B2(n5920), .C1(n47), .C2(n5930), .A(n5243), 
        .ZN(n5238) );
  AOI22_X1 U1836 ( .A1(n5934), .A2(n2613), .B1(n5942), .B2(n2614), .ZN(n5243)
         );
  OAI221_X1 U1837 ( .B1(n2005), .B2(n6051), .C1(n44), .C2(n6058), .A(n5235), 
        .ZN(n5230) );
  AOI22_X1 U1838 ( .A1(n6062), .A2(n2597), .B1(n6071), .B2(n2598), .ZN(n5235)
         );
  OAI221_X1 U1839 ( .B1(n2304), .B2(n5919), .C1(n40), .C2(n5931), .A(n5225), 
        .ZN(n5220) );
  AOI22_X1 U1840 ( .A1(n5938), .A2(n2579), .B1(n5943), .B2(n2580), .ZN(n5225)
         );
  OAI221_X1 U1841 ( .B1(n2285), .B2(n5922), .C1(n96), .C2(n5930), .A(n5369), 
        .ZN(n5364) );
  AOI22_X1 U1842 ( .A1(n5939), .A2(n4452), .B1(n5947), .B2(n4453), .ZN(n5369)
         );
  OAI221_X1 U1843 ( .B1(n1984), .B2(n6049), .C1(n93), .C2(n6056), .A(n5361), 
        .ZN(n5356) );
  AOI22_X1 U1844 ( .A1(n6067), .A2(n4436), .B1(n6073), .B2(n4437), .ZN(n5361)
         );
  OAI221_X1 U1845 ( .B1(n2284), .B2(n5923), .C1(n89), .C2(n5929), .A(n5351), 
        .ZN(n5346) );
  AOI22_X1 U1846 ( .A1(n5938), .A2(n4418), .B1(n5947), .B2(n4419), .ZN(n5351)
         );
  OAI221_X1 U1847 ( .B1(n1983), .B2(n6050), .C1(n86), .C2(n6057), .A(n5343), 
        .ZN(n5338) );
  AOI22_X1 U1848 ( .A1(n6066), .A2(n4402), .B1(n6075), .B2(n4403), .ZN(n5343)
         );
  OAI221_X1 U1849 ( .B1(n2283), .B2(n5922), .C1(n82), .C2(n5930), .A(n5333), 
        .ZN(n5328) );
  AOI22_X1 U1850 ( .A1(n5937), .A2(n4384), .B1(n5942), .B2(n4385), .ZN(n5333)
         );
  OAI221_X1 U1851 ( .B1(n1982), .B2(n6051), .C1(n79), .C2(n6056), .A(n5325), 
        .ZN(n5320) );
  AOI22_X1 U1852 ( .A1(n6065), .A2(n4368), .B1(n6075), .B2(n4369), .ZN(n5325)
         );
  OAI221_X1 U1853 ( .B1(n2282), .B2(n5922), .C1(n75), .C2(n5930), .A(n5315), 
        .ZN(n5310) );
  AOI22_X1 U1854 ( .A1(n5936), .A2(n4350), .B1(n5943), .B2(n4351), .ZN(n5315)
         );
  OAI221_X1 U1855 ( .B1(n1981), .B2(n6049), .C1(n72), .C2(n6057), .A(n5307), 
        .ZN(n5302) );
  AOI22_X1 U1856 ( .A1(n6064), .A2(n4334), .B1(n6075), .B2(n4335), .ZN(n5307)
         );
  OAI221_X1 U1857 ( .B1(n2306), .B2(n5921), .C1(n68), .C2(n5931), .A(n5297), 
        .ZN(n5292) );
  AOI22_X1 U1858 ( .A1(n5933), .A2(n4316), .B1(n5941), .B2(n4317), .ZN(n5297)
         );
  OAI221_X1 U1859 ( .B1(n2006), .B2(n6049), .C1(n65), .C2(n6059), .A(n5289), 
        .ZN(n5284) );
  AOI22_X1 U1860 ( .A1(n6061), .A2(n4300), .B1(n6070), .B2(n4301), .ZN(n5289)
         );
  OAI221_X1 U1861 ( .B1(n2281), .B2(n5923), .C1(n61), .C2(n5931), .A(n5279), 
        .ZN(n5274) );
  AOI22_X1 U1862 ( .A1(n5938), .A2(n3706), .B1(n5947), .B2(n3707), .ZN(n5279)
         );
  OAI221_X1 U1863 ( .B1(n1980), .B2(n6050), .C1(n58), .C2(n6059), .A(n5271), 
        .ZN(n5266) );
  AOI22_X1 U1864 ( .A1(n6066), .A2(n3690), .B1(n6073), .B2(n3691), .ZN(n5271)
         );
  OAI221_X1 U1865 ( .B1(n1925), .B2(n6018), .C1(n8), .C2(n6023), .A(n5146), 
        .ZN(n5139) );
  AOI22_X1 U1866 ( .A1(n6032), .A2(n2430), .B1(n6041), .B2(n2431), .ZN(n5146)
         );
  OAI221_X1 U1867 ( .B1(n1881), .B2(n6018), .C1(n50), .C2(n6027), .A(n5254), 
        .ZN(n5247) );
  AOI22_X1 U1868 ( .A1(n6030), .A2(n2634), .B1(n6037), .B2(n2635), .ZN(n5254)
         );
  OAI221_X1 U1869 ( .B1(n1935), .B2(n6018), .C1(n43), .C2(n6027), .A(n5236), 
        .ZN(n5229) );
  AOI22_X1 U1870 ( .A1(n6031), .A2(n2600), .B1(n6039), .B2(n2601), .ZN(n5236)
         );
  OAI221_X1 U1871 ( .B1(n1893), .B2(n6016), .C1(n99), .C2(n6026), .A(n5380), 
        .ZN(n5373) );
  AOI22_X1 U1872 ( .A1(n6035), .A2(n4473), .B1(n6041), .B2(n4474), .ZN(n5380)
         );
  OAI221_X1 U1873 ( .B1(n1937), .B2(n6019), .C1(n64), .C2(n6026), .A(n5290), 
        .ZN(n5283) );
  AOI22_X1 U1874 ( .A1(n6030), .A2(n4303), .B1(n6037), .B2(n4304), .ZN(n5290)
         );
  OAI221_X1 U1875 ( .B1(n1883), .B2(n6019), .C1(n57), .C2(n6025), .A(n5272), 
        .ZN(n5265) );
  AOI22_X1 U1876 ( .A1(n6034), .A2(n3693), .B1(n6043), .B2(n3694), .ZN(n5272)
         );
  INV_X1 U1877 ( .A(ADD_RD1[4]), .ZN(n5705) );
  INV_X1 U1878 ( .A(RD1), .ZN(n5710) );
  INV_X1 U1879 ( .A(ADD_RD1[0]), .ZN(n5691) );
  INV_X1 U1880 ( .A(ADD_RD1[3]), .ZN(n5692) );
  NAND2_X1 U1881 ( .A1(n5677), .A2(n5678), .ZN(OUT1[0]) );
  NOR4_X1 U1882 ( .A1(n5679), .A2(n5680), .A3(n5681), .A4(n5682), .ZN(n5678)
         );
  NOR4_X1 U1883 ( .A1(n5697), .A2(n5698), .A3(n5699), .A4(n5700), .ZN(n5677)
         );
  OAI221_X1 U1884 ( .B1(n444), .B2(n6079), .C1(n2094), .C2(n6089), .A(n5688), 
        .ZN(n5681) );
  NAND2_X1 U1885 ( .A1(n5245), .A2(n5246), .ZN(OUT1[31]) );
  NOR4_X1 U1886 ( .A1(n5247), .A2(n5248), .A3(n5249), .A4(n5250), .ZN(n5246)
         );
  NOR4_X1 U1887 ( .A1(n5255), .A2(n5256), .A3(n5257), .A4(n5258), .ZN(n5245)
         );
  OAI221_X1 U1888 ( .B1(n2040), .B2(n6083), .C1(n52), .C2(n6090), .A(n5252), 
        .ZN(n5249) );
  NAND2_X1 U1889 ( .A1(n5317), .A2(n5318), .ZN(OUT1[28]) );
  NOR4_X1 U1890 ( .A1(n5319), .A2(n5320), .A3(n5321), .A4(n5322), .ZN(n5318)
         );
  NOR4_X1 U1891 ( .A1(n5327), .A2(n5328), .A3(n5329), .A4(n5330), .ZN(n5317)
         );
  OAI221_X1 U1892 ( .B1(n1887), .B2(n6017), .C1(n78), .C2(n6026), .A(n5326), 
        .ZN(n5319) );
  NAND2_X1 U1893 ( .A1(n5659), .A2(n5660), .ZN(OUT1[10]) );
  NOR4_X1 U1894 ( .A1(n5661), .A2(n5662), .A3(n5663), .A4(n5664), .ZN(n5660)
         );
  NOR4_X1 U1895 ( .A1(n5669), .A2(n5670), .A3(n5671), .A4(n5672), .ZN(n5659)
         );
  OAI221_X1 U1896 ( .B1(n437), .B2(n6080), .C1(n2086), .C2(n6086), .A(n5666), 
        .ZN(n5663) );
  NAND2_X1 U1897 ( .A1(n5227), .A2(n5228), .ZN(OUT1[3]) );
  NOR4_X1 U1898 ( .A1(n5229), .A2(n5230), .A3(n5231), .A4(n5232), .ZN(n5228)
         );
  NOR4_X1 U1899 ( .A1(n5237), .A2(n5238), .A3(n5239), .A4(n5240), .ZN(n5227)
         );
  OAI221_X1 U1900 ( .B1(n2065), .B2(n6083), .C1(n45), .C2(n6087), .A(n5234), 
        .ZN(n5231) );
  NAND2_X1 U1901 ( .A1(n5299), .A2(n5300), .ZN(OUT1[29]) );
  NOR4_X1 U1902 ( .A1(n5301), .A2(n5302), .A3(n5303), .A4(n5304), .ZN(n5300)
         );
  NOR4_X1 U1903 ( .A1(n5309), .A2(n5310), .A3(n5311), .A4(n5312), .ZN(n5299)
         );
  OAI221_X1 U1904 ( .B1(n1885), .B2(n6017), .C1(n71), .C2(n6026), .A(n5308), 
        .ZN(n5301) );
  NAND2_X1 U1905 ( .A1(n5641), .A2(n5642), .ZN(OUT1[11]) );
  NOR4_X1 U1906 ( .A1(n5643), .A2(n5644), .A3(n5645), .A4(n5646), .ZN(n5642)
         );
  NOR4_X1 U1907 ( .A1(n5651), .A2(n5652), .A3(n5653), .A4(n5654), .ZN(n5641)
         );
  OAI221_X1 U1908 ( .B1(n430), .B2(n6078), .C1(n2085), .C2(n6087), .A(n5648), 
        .ZN(n5645) );
  NAND2_X1 U1909 ( .A1(n5353), .A2(n5354), .ZN(OUT1[26]) );
  NOR4_X1 U1910 ( .A1(n5355), .A2(n5356), .A3(n5357), .A4(n5358), .ZN(n5354)
         );
  NOR4_X1 U1911 ( .A1(n5363), .A2(n5364), .A3(n5365), .A4(n5366), .ZN(n5353)
         );
  OAI221_X1 U1912 ( .B1(n1891), .B2(n6017), .C1(n92), .C2(n6025), .A(n5362), 
        .ZN(n5355) );
  NAND2_X1 U1913 ( .A1(n5281), .A2(n5282), .ZN(OUT1[2]) );
  NOR4_X1 U1914 ( .A1(n5283), .A2(n5284), .A3(n5285), .A4(n5286), .ZN(n5282)
         );
  NOR4_X1 U1915 ( .A1(n5291), .A2(n5292), .A3(n5293), .A4(n5294), .ZN(n5281)
         );
  OAI221_X1 U1916 ( .B1(n2066), .B2(n6082), .C1(n66), .C2(n6091), .A(n5288), 
        .ZN(n5285) );
  NAND2_X1 U1917 ( .A1(n5335), .A2(n5336), .ZN(OUT1[27]) );
  NOR4_X1 U1918 ( .A1(n5337), .A2(n5338), .A3(n5339), .A4(n5340), .ZN(n5336)
         );
  NOR4_X1 U1919 ( .A1(n5345), .A2(n5346), .A3(n5347), .A4(n5348), .ZN(n5335)
         );
  OAI221_X1 U1920 ( .B1(n1889), .B2(n6019), .C1(n85), .C2(n6025), .A(n5344), 
        .ZN(n5337) );
  NAND2_X1 U1921 ( .A1(n5263), .A2(n5264), .ZN(OUT1[30]) );
  NOR4_X1 U1922 ( .A1(n5265), .A2(n5266), .A3(n5267), .A4(n5268), .ZN(n5264)
         );
  NOR4_X1 U1923 ( .A1(n5273), .A2(n5274), .A3(n5275), .A4(n5276), .ZN(n5263)
         );
  OAI221_X1 U1924 ( .B1(n2041), .B2(n6080), .C1(n59), .C2(n6091), .A(n5270), 
        .ZN(n5267) );
  INV_X1 U1925 ( .A(ADD_RD1[1]), .ZN(n5709) );
  INV_X1 U1926 ( .A(ADD_RD1[2]), .ZN(n5712) );
  NOR3_X1 U1927 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n5059) );
  NOR3_X1 U1928 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n5053), .ZN(n5058) );
  NOR3_X1 U1929 ( .A1(n5053), .A2(ADD_RD2[3]), .A3(n5075), .ZN(n5071) );
  NOR3_X1 U1930 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n5075), .ZN(n5070) );
  NOR3_X1 U1931 ( .A1(n5054), .A2(ADD_RD2[0]), .A3(n5075), .ZN(n5079) );
  NAND2_X1 U1932 ( .A1(ADD_WR[1]), .A2(n2341), .ZN(n1970) );
  OAI221_X1 U1933 ( .B1(n445), .B2(n6330), .C1(n2153), .C2(n6338), .A(n5041), 
        .ZN(n5040) );
  AOI22_X1 U1934 ( .A1(n6344), .A2(n5042), .B1(n6346), .B2(n5043), .ZN(n5041)
         );
  OAI221_X1 U1935 ( .B1(n448), .B2(n6214), .C1(n2242), .C2(n6222), .A(n5067), 
        .ZN(n5066) );
  AOI22_X1 U1936 ( .A1(n6233), .A2(n5068), .B1(n6237), .B2(n5069), .ZN(n5067)
         );
  OAI221_X1 U1937 ( .B1(n438), .B2(n6329), .C1(n2147), .C2(n6339), .A(n5007), 
        .ZN(n5006) );
  AOI22_X1 U1938 ( .A1(n6345), .A2(n5008), .B1(n6347), .B2(n5009), .ZN(n5007)
         );
  OAI221_X1 U1939 ( .B1(n441), .B2(n6213), .C1(n2236), .C2(n6223), .A(n5023), 
        .ZN(n5022) );
  AOI22_X1 U1940 ( .A1(n6232), .A2(n5024), .B1(n6240), .B2(n5025), .ZN(n5023)
         );
  OAI221_X1 U1941 ( .B1(n431), .B2(n6334), .C1(n2146), .C2(n6341), .A(n4973), 
        .ZN(n4972) );
  AOI22_X1 U1942 ( .A1(n2357), .A2(n4974), .B1(n2359), .B2(n4975), .ZN(n4973)
         );
  OAI221_X1 U1943 ( .B1(n434), .B2(n6218), .C1(n2235), .C2(n6225), .A(n4989), 
        .ZN(n4988) );
  AOI22_X1 U1944 ( .A1(n6229), .A2(n4990), .B1(n6237), .B2(n4991), .ZN(n4989)
         );
  OAI221_X1 U1945 ( .B1(n424), .B2(n6333), .C1(n2145), .C2(n6342), .A(n4939), 
        .ZN(n4938) );
  AOI22_X1 U1946 ( .A1(n6344), .A2(n4940), .B1(n6346), .B2(n4941), .ZN(n4939)
         );
  OAI221_X1 U1947 ( .B1(n427), .B2(n6217), .C1(n2234), .C2(n6226), .A(n4955), 
        .ZN(n4954) );
  AOI22_X1 U1948 ( .A1(n6229), .A2(n4956), .B1(n6237), .B2(n4957), .ZN(n4955)
         );
  OAI221_X1 U1949 ( .B1(n2127), .B2(n6333), .C1(n67), .C2(n6341), .A(n3717), 
        .ZN(n3716) );
  AOI22_X1 U1950 ( .A1(n6345), .A2(n3718), .B1(n6347), .B2(n3719), .ZN(n3717)
         );
  OAI221_X1 U1951 ( .B1(n2272), .B2(n6217), .C1(n70), .C2(n6225), .A(n4309), 
        .ZN(n4308) );
  AOI22_X1 U1952 ( .A1(n6233), .A2(n4310), .B1(n6237), .B2(n4311), .ZN(n4309)
         );
  OAI221_X1 U1953 ( .B1(n2126), .B2(n6334), .C1(n46), .C2(n6343), .A(n2590), 
        .ZN(n2589) );
  AOI22_X1 U1954 ( .A1(n6345), .A2(n2591), .B1(n6347), .B2(n2592), .ZN(n2590)
         );
  OAI221_X1 U1955 ( .B1(n2271), .B2(n6218), .C1(n49), .C2(n6227), .A(n2606), 
        .ZN(n2605) );
  AOI22_X1 U1956 ( .A1(n6229), .A2(n2607), .B1(n6237), .B2(n2608), .ZN(n2606)
         );
  OAI221_X1 U1957 ( .B1(n2125), .B2(n6334), .C1(n39), .C2(n6342), .A(n2556), 
        .ZN(n2555) );
  AOI22_X1 U1958 ( .A1(n2357), .A2(n2557), .B1(n2359), .B2(n2558), .ZN(n2556)
         );
  OAI221_X1 U1959 ( .B1(n2270), .B2(n6218), .C1(n42), .C2(n6226), .A(n2572), 
        .ZN(n2571) );
  AOI22_X1 U1960 ( .A1(n6229), .A2(n2573), .B1(n6238), .B2(n2574), .ZN(n2572)
         );
  OAI221_X1 U1961 ( .B1(n2120), .B2(n6331), .C1(n4), .C2(n6340), .A(n2356), 
        .ZN(n2353) );
  AOI22_X1 U1962 ( .A1(n6345), .A2(n2358), .B1(n6347), .B2(n2360), .ZN(n2356)
         );
  OAI221_X1 U1963 ( .B1(n2265), .B2(n6215), .C1(n7), .C2(n6224), .A(n2388), 
        .ZN(n2385) );
  AOI22_X1 U1964 ( .A1(n6232), .A2(n2390), .B1(n6241), .B2(n2392), .ZN(n2388)
         );
  OAI221_X1 U1965 ( .B1(n2106), .B2(n6333), .C1(n95), .C2(n6340), .A(n4429), 
        .ZN(n4428) );
  AOI22_X1 U1966 ( .A1(n6344), .A2(n4430), .B1(n6346), .B2(n4431), .ZN(n4429)
         );
  OAI221_X1 U1967 ( .B1(n2251), .B2(n6217), .C1(n98), .C2(n6224), .A(n4445), 
        .ZN(n4444) );
  AOI22_X1 U1968 ( .A1(n6235), .A2(n4446), .B1(n6243), .B2(n4447), .ZN(n4445)
         );
  OAI221_X1 U1969 ( .B1(n2105), .B2(n6333), .C1(n88), .C2(n6340), .A(n4395), 
        .ZN(n4394) );
  AOI22_X1 U1970 ( .A1(n6345), .A2(n4396), .B1(n6347), .B2(n4397), .ZN(n4395)
         );
  OAI221_X1 U1971 ( .B1(n2250), .B2(n6217), .C1(n91), .C2(n6224), .A(n4411), 
        .ZN(n4410) );
  AOI22_X1 U1972 ( .A1(n6235), .A2(n4412), .B1(n6243), .B2(n4413), .ZN(n4411)
         );
  OAI221_X1 U1973 ( .B1(n2104), .B2(n6333), .C1(n81), .C2(n6341), .A(n4361), 
        .ZN(n4360) );
  AOI22_X1 U1974 ( .A1(n2357), .A2(n4362), .B1(n2359), .B2(n4363), .ZN(n4361)
         );
  OAI221_X1 U1975 ( .B1(n2249), .B2(n6217), .C1(n84), .C2(n6225), .A(n4377), 
        .ZN(n4376) );
  AOI22_X1 U1976 ( .A1(n6235), .A2(n4378), .B1(n6243), .B2(n4379), .ZN(n4377)
         );
  OAI221_X1 U1977 ( .B1(n2103), .B2(n6334), .C1(n74), .C2(n6342), .A(n4327), 
        .ZN(n4326) );
  AOI22_X1 U1978 ( .A1(n6344), .A2(n4328), .B1(n6346), .B2(n4329), .ZN(n4327)
         );
  OAI221_X1 U1979 ( .B1(n2248), .B2(n6218), .C1(n77), .C2(n6226), .A(n4343), 
        .ZN(n4342) );
  AOI22_X1 U1980 ( .A1(n6235), .A2(n4344), .B1(n6243), .B2(n4345), .ZN(n4343)
         );
  OAI221_X1 U1981 ( .B1(n2102), .B2(n6335), .C1(n60), .C2(n6342), .A(n3683), 
        .ZN(n3682) );
  AOI22_X1 U1982 ( .A1(n2357), .A2(n3684), .B1(n2359), .B2(n3685), .ZN(n3683)
         );
  OAI221_X1 U1983 ( .B1(n2247), .B2(n6219), .C1(n63), .C2(n6226), .A(n3699), 
        .ZN(n3698) );
  AOI22_X1 U1984 ( .A1(n6229), .A2(n3700), .B1(n6240), .B2(n3701), .ZN(n3699)
         );
  OAI221_X1 U1985 ( .B1(n2101), .B2(n6335), .C1(n53), .C2(n6343), .A(n2624), 
        .ZN(n2623) );
  AOI22_X1 U1986 ( .A1(n6344), .A2(n2625), .B1(n6346), .B2(n2626), .ZN(n2624)
         );
  OAI221_X1 U1987 ( .B1(n2246), .B2(n6219), .C1(n56), .C2(n6227), .A(n2640), 
        .ZN(n2639) );
  AOI22_X1 U1988 ( .A1(n6230), .A2(n2641), .B1(n6239), .B2(n2642), .ZN(n2640)
         );
  OAI221_X1 U1989 ( .B1(n444), .B2(n6310), .C1(n2094), .C2(n6318), .A(n5048), 
        .ZN(n5039) );
  AOI22_X1 U1990 ( .A1(n6324), .A2(n5049), .B1(n6326), .B2(n5050), .ZN(n5048)
         );
  OAI221_X1 U1991 ( .B1(n447), .B2(n6182), .C1(n2182), .C2(n6190), .A(n5072), 
        .ZN(n5065) );
  AOI22_X1 U1992 ( .A1(n6201), .A2(n5073), .B1(n6205), .B2(n5074), .ZN(n5072)
         );
  OAI221_X1 U1993 ( .B1(n437), .B2(n6309), .C1(n2086), .C2(n6319), .A(n5010), 
        .ZN(n5005) );
  AOI22_X1 U1994 ( .A1(n6325), .A2(n5011), .B1(n6327), .B2(n5012), .ZN(n5010)
         );
  OAI221_X1 U1995 ( .B1(n440), .B2(n6181), .C1(n2176), .C2(n6191), .A(n5026), 
        .ZN(n5021) );
  AOI22_X1 U1996 ( .A1(n6200), .A2(n5027), .B1(n6207), .B2(n5028), .ZN(n5026)
         );
  OAI221_X1 U1997 ( .B1(n430), .B2(n6313), .C1(n2085), .C2(n6321), .A(n4976), 
        .ZN(n4971) );
  AOI22_X1 U1998 ( .A1(n2364), .A2(n4977), .B1(n2366), .B2(n4978), .ZN(n4976)
         );
  OAI221_X1 U1999 ( .B1(n433), .B2(n6186), .C1(n2175), .C2(n6193), .A(n4992), 
        .ZN(n4987) );
  AOI22_X1 U2000 ( .A1(n6197), .A2(n4993), .B1(n6205), .B2(n4994), .ZN(n4992)
         );
  OAI221_X1 U2001 ( .B1(n423), .B2(n6314), .C1(n2084), .C2(n6322), .A(n4942), 
        .ZN(n4937) );
  AOI22_X1 U2002 ( .A1(n6324), .A2(n4943), .B1(n6326), .B2(n4944), .ZN(n4942)
         );
  OAI221_X1 U2003 ( .B1(n426), .B2(n6185), .C1(n2174), .C2(n6194), .A(n4958), 
        .ZN(n4953) );
  AOI22_X1 U2004 ( .A1(n6197), .A2(n4959), .B1(n6205), .B2(n4960), .ZN(n4958)
         );
  OAI221_X1 U2005 ( .B1(n2066), .B2(n6313), .C1(n66), .C2(n6321), .A(n3720), 
        .ZN(n3715) );
  AOI22_X1 U2006 ( .A1(n6325), .A2(n3721), .B1(n6327), .B2(n4298), .ZN(n3720)
         );
  OAI221_X1 U2007 ( .B1(n2212), .B2(n6185), .C1(n69), .C2(n6193), .A(n4312), 
        .ZN(n4307) );
  AOI22_X1 U2008 ( .A1(n6201), .A2(n4313), .B1(n6205), .B2(n4314), .ZN(n4312)
         );
  OAI221_X1 U2009 ( .B1(n2065), .B2(n6314), .C1(n45), .C2(n6323), .A(n2593), 
        .ZN(n2588) );
  AOI22_X1 U2010 ( .A1(n6325), .A2(n2594), .B1(n6327), .B2(n2595), .ZN(n2593)
         );
  OAI221_X1 U2011 ( .B1(n2211), .B2(n6186), .C1(n48), .C2(n6195), .A(n2609), 
        .ZN(n2604) );
  AOI22_X1 U2012 ( .A1(n6197), .A2(n2610), .B1(n6205), .B2(n2611), .ZN(n2609)
         );
  OAI221_X1 U2013 ( .B1(n2210), .B2(n6186), .C1(n41), .C2(n6194), .A(n2575), 
        .ZN(n2570) );
  AOI22_X1 U2014 ( .A1(n6197), .A2(n2576), .B1(n6206), .B2(n2577), .ZN(n2575)
         );
  OAI221_X1 U2015 ( .B1(n2205), .B2(n6183), .C1(n6), .C2(n6192), .A(n2395), 
        .ZN(n2384) );
  AOI22_X1 U2016 ( .A1(n6200), .A2(n2397), .B1(n6209), .B2(n2399), .ZN(n2395)
         );
  OAI221_X1 U2017 ( .B1(n2045), .B2(n6313), .C1(n94), .C2(n6320), .A(n4432), 
        .ZN(n4427) );
  AOI22_X1 U2018 ( .A1(n6324), .A2(n4433), .B1(n6326), .B2(n4434), .ZN(n4432)
         );
  OAI221_X1 U2019 ( .B1(n2191), .B2(n6185), .C1(n97), .C2(n6192), .A(n4448), 
        .ZN(n4443) );
  AOI22_X1 U2020 ( .A1(n6203), .A2(n4449), .B1(n6211), .B2(n4450), .ZN(n4448)
         );
  OAI221_X1 U2021 ( .B1(n2044), .B2(n6311), .C1(n87), .C2(n6320), .A(n4398), 
        .ZN(n4393) );
  AOI22_X1 U2022 ( .A1(n6325), .A2(n4399), .B1(n6327), .B2(n4400), .ZN(n4398)
         );
  OAI221_X1 U2023 ( .B1(n2190), .B2(n6185), .C1(n90), .C2(n6192), .A(n4414), 
        .ZN(n4409) );
  AOI22_X1 U2024 ( .A1(n6203), .A2(n4415), .B1(n6211), .B2(n4416), .ZN(n4414)
         );
  OAI221_X1 U2025 ( .B1(n2043), .B2(n6315), .C1(n80), .C2(n6321), .A(n4364), 
        .ZN(n4359) );
  AOI22_X1 U2026 ( .A1(n2364), .A2(n4365), .B1(n2366), .B2(n4366), .ZN(n4364)
         );
  OAI221_X1 U2027 ( .B1(n2189), .B2(n6185), .C1(n83), .C2(n6193), .A(n4380), 
        .ZN(n4375) );
  AOI22_X1 U2028 ( .A1(n6203), .A2(n4381), .B1(n6211), .B2(n4382), .ZN(n4380)
         );
  OAI221_X1 U2029 ( .B1(n2042), .B2(n6315), .C1(n73), .C2(n6322), .A(n4330), 
        .ZN(n4325) );
  AOI22_X1 U2030 ( .A1(n6324), .A2(n4331), .B1(n6326), .B2(n4332), .ZN(n4330)
         );
  OAI221_X1 U2031 ( .B1(n2188), .B2(n6186), .C1(n76), .C2(n6194), .A(n4346), 
        .ZN(n4341) );
  AOI22_X1 U2032 ( .A1(n6203), .A2(n4347), .B1(n6211), .B2(n4348), .ZN(n4346)
         );
  OAI221_X1 U2033 ( .B1(n2041), .B2(n6315), .C1(n59), .C2(n6322), .A(n3686), 
        .ZN(n2656) );
  AOI22_X1 U2034 ( .A1(n2364), .A2(n3687), .B1(n2366), .B2(n3688), .ZN(n3686)
         );
  OAI221_X1 U2035 ( .B1(n2187), .B2(n6187), .C1(n62), .C2(n6194), .A(n3702), 
        .ZN(n3697) );
  AOI22_X1 U2036 ( .A1(n6197), .A2(n3703), .B1(n6208), .B2(n3704), .ZN(n3702)
         );
  OAI221_X1 U2037 ( .B1(n2040), .B2(n6314), .C1(n52), .C2(n6323), .A(n2627), 
        .ZN(n2622) );
  AOI22_X1 U2038 ( .A1(n6324), .A2(n2628), .B1(n6326), .B2(n2629), .ZN(n2627)
         );
  OAI221_X1 U2039 ( .B1(n2186), .B2(n6187), .C1(n55), .C2(n6195), .A(n2643), 
        .ZN(n2638) );
  AOI22_X1 U2040 ( .A1(n6198), .A2(n2644), .B1(n6207), .B2(n2645), .ZN(n2643)
         );
  OAI221_X1 U2041 ( .B1(n443), .B2(n6278), .C1(n2033), .C2(n6286), .A(n5055), 
        .ZN(n5038) );
  AOI22_X1 U2042 ( .A1(n6293), .A2(n5056), .B1(n6302), .B2(n5057), .ZN(n5055)
         );
  OAI221_X1 U2043 ( .B1(n446), .B2(n6150), .C1(n2332), .C2(n6158), .A(n5076), 
        .ZN(n5064) );
  AOI22_X1 U2044 ( .A1(n6169), .A2(n5077), .B1(n6173), .B2(n5078), .ZN(n5076)
         );
  OAI221_X1 U2045 ( .B1(n436), .B2(n6280), .C1(n2026), .C2(n6289), .A(n5013), 
        .ZN(n5004) );
  AOI22_X1 U2046 ( .A1(n6293), .A2(n5014), .B1(n6304), .B2(n5015), .ZN(n5013)
         );
  OAI221_X1 U2047 ( .B1(n439), .B2(n6149), .C1(n2326), .C2(n6159), .A(n5029), 
        .ZN(n5020) );
  AOI22_X1 U2048 ( .A1(n6168), .A2(n5030), .B1(n6176), .B2(n5031), .ZN(n5029)
         );
  OAI221_X1 U2049 ( .B1(n429), .B2(n6281), .C1(n2025), .C2(n6288), .A(n4979), 
        .ZN(n4970) );
  AOI22_X1 U2050 ( .A1(n6299), .A2(n4980), .B1(n6301), .B2(n4981), .ZN(n4979)
         );
  OAI221_X1 U2051 ( .B1(n432), .B2(n6154), .C1(n2325), .C2(n6161), .A(n4995), 
        .ZN(n4986) );
  AOI22_X1 U2052 ( .A1(n6165), .A2(n4996), .B1(n6173), .B2(n4997), .ZN(n4995)
         );
  OAI221_X1 U2053 ( .B1(n425), .B2(n6153), .C1(n2324), .C2(n6162), .A(n4961), 
        .ZN(n4952) );
  AOI22_X1 U2054 ( .A1(n6165), .A2(n4962), .B1(n6173), .B2(n4963), .ZN(n4961)
         );
  OAI221_X1 U2055 ( .B1(n442), .B2(n6247), .C1(n1966), .C2(n6253), .A(n5060), 
        .ZN(n5037) );
  AOI22_X1 U2056 ( .A1(n6261), .A2(n5061), .B1(n6270), .B2(n5062), .ZN(n5060)
         );
  OAI221_X1 U2057 ( .B1(n4295), .B2(n6117), .C1(n4294), .C2(n6127), .A(n5083), 
        .ZN(n5063) );
  AOI22_X1 U2058 ( .A1(n6133), .A2(n5084), .B1(n6141), .B2(n5085), .ZN(n5083)
         );
  OAI221_X1 U2059 ( .B1(n4097), .B2(n6119), .C1(n4096), .C2(n6129), .A(n4692), 
        .ZN(n4679) );
  AOI22_X1 U2060 ( .A1(n6137), .A2(n4693), .B1(n6142), .B2(n4694), .ZN(n4692)
         );
  OAI221_X1 U2061 ( .B1(n3899), .B2(n6121), .C1(n3898), .C2(n6129), .A(n4318), 
        .ZN(n4305) );
  AOI22_X1 U2062 ( .A1(n6133), .A2(n4319), .B1(n6141), .B2(n4320), .ZN(n4318)
         );
  OAI221_X1 U2063 ( .B1(n3845), .B2(n6122), .C1(n3844), .C2(n6131), .A(n2615), 
        .ZN(n2602) );
  AOI22_X1 U2064 ( .A1(n6134), .A2(n2616), .B1(n6145), .B2(n2617), .ZN(n2615)
         );
  OAI221_X1 U2065 ( .B1(n3827), .B2(n6123), .C1(n3826), .C2(n6130), .A(n2581), 
        .ZN(n2568) );
  AOI22_X1 U2066 ( .A1(n6134), .A2(n2582), .B1(n6142), .B2(n2583), .ZN(n2581)
         );
  OAI221_X1 U2067 ( .B1(n3809), .B2(n6123), .C1(n3808), .C2(n6131), .A(n2547), 
        .ZN(n2534) );
  AOI22_X1 U2068 ( .A1(n6133), .A2(n2548), .B1(n6142), .B2(n2549), .ZN(n2547)
         );
  OAI221_X1 U2069 ( .B1(n3791), .B2(n6117), .C1(n3790), .C2(n6127), .A(n2513), 
        .ZN(n2500) );
  AOI22_X1 U2070 ( .A1(n6135), .A2(n2514), .B1(n6143), .B2(n2515), .ZN(n2513)
         );
  OAI221_X1 U2071 ( .B1(n3773), .B2(n6117), .C1(n3772), .C2(n6128), .A(n2479), 
        .ZN(n2466) );
  AOI22_X1 U2072 ( .A1(n6134), .A2(n2480), .B1(n6144), .B2(n2481), .ZN(n2479)
         );
  OAI221_X1 U2073 ( .B1(n3755), .B2(n6118), .C1(n3754), .C2(n6126), .A(n2445), 
        .ZN(n2432) );
  AOI22_X1 U2074 ( .A1(n6136), .A2(n2446), .B1(n6143), .B2(n2447), .ZN(n2445)
         );
  OAI221_X1 U2075 ( .B1(n3737), .B2(n6120), .C1(n3736), .C2(n6131), .A(n2409), 
        .ZN(n2382) );
  AOI22_X1 U2076 ( .A1(n6137), .A2(n2411), .B1(n6145), .B2(n2413), .ZN(n2409)
         );
  OAI221_X1 U2077 ( .B1(n435), .B2(n6249), .C1(n1959), .C2(n6259), .A(n5016), 
        .ZN(n5003) );
  AOI22_X1 U2078 ( .A1(n6261), .A2(n5017), .B1(n6272), .B2(n5018), .ZN(n5016)
         );
  OAI221_X1 U2079 ( .B1(n4277), .B2(n6118), .C1(n4276), .C2(n6128), .A(n5032), 
        .ZN(n5019) );
  AOI22_X1 U2080 ( .A1(n6133), .A2(n5033), .B1(n6144), .B2(n5034), .ZN(n5032)
         );
  OAI221_X1 U2081 ( .B1(n428), .B2(n6248), .C1(n1958), .C2(n6255), .A(n4982), 
        .ZN(n4969) );
  AOI22_X1 U2082 ( .A1(n6264), .A2(n4983), .B1(n6269), .B2(n4984), .ZN(n4982)
         );
  OAI221_X1 U2083 ( .B1(n4259), .B2(n6118), .C1(n4258), .C2(n6129), .A(n4998), 
        .ZN(n4985) );
  AOI22_X1 U2084 ( .A1(n6136), .A2(n4999), .B1(n6141), .B2(n5000), .ZN(n4998)
         );
  OAI221_X1 U2085 ( .B1(n4241), .B2(n6119), .C1(n4240), .C2(n6130), .A(n4964), 
        .ZN(n4951) );
  AOI22_X1 U2086 ( .A1(n6134), .A2(n4965), .B1(n6141), .B2(n4966), .ZN(n4964)
         );
  OAI221_X1 U2087 ( .B1(n4223), .B2(n6123), .C1(n4222), .C2(n6127), .A(n4930), 
        .ZN(n4917) );
  AOI22_X1 U2088 ( .A1(n6134), .A2(n4931), .B1(n6142), .B2(n4932), .ZN(n4930)
         );
  OAI221_X1 U2089 ( .B1(n4205), .B2(n6119), .C1(n4204), .C2(n6126), .A(n4896), 
        .ZN(n4883) );
  AOI22_X1 U2090 ( .A1(n6137), .A2(n4897), .B1(n6142), .B2(n4898), .ZN(n4896)
         );
  OAI221_X1 U2091 ( .B1(n4187), .B2(n6120), .C1(n4186), .C2(n6127), .A(n4862), 
        .ZN(n4849) );
  AOI22_X1 U2092 ( .A1(n6135), .A2(n4863), .B1(n6143), .B2(n4864), .ZN(n4862)
         );
  OAI221_X1 U2093 ( .B1(n4169), .B2(n6120), .C1(n4168), .C2(n6127), .A(n4828), 
        .ZN(n4815) );
  AOI22_X1 U2094 ( .A1(n6136), .A2(n4829), .B1(n6144), .B2(n4830), .ZN(n4828)
         );
  OAI221_X1 U2095 ( .B1(n4151), .B2(n6121), .C1(n4150), .C2(n6128), .A(n4794), 
        .ZN(n4781) );
  AOI22_X1 U2096 ( .A1(n6136), .A2(n4795), .B1(n6144), .B2(n4796), .ZN(n4794)
         );
  OAI221_X1 U2097 ( .B1(n4133), .B2(n6121), .C1(n4132), .C2(n6129), .A(n4760), 
        .ZN(n4747) );
  AOI22_X1 U2098 ( .A1(n6135), .A2(n4761), .B1(n6145), .B2(n4762), .ZN(n4760)
         );
  OAI221_X1 U2099 ( .B1(n4115), .B2(n6119), .C1(n4114), .C2(n6128), .A(n4726), 
        .ZN(n4713) );
  AOI22_X1 U2100 ( .A1(n6137), .A2(n4727), .B1(n6145), .B2(n4728), .ZN(n4726)
         );
  OAI221_X1 U2101 ( .B1(n4079), .B2(n6121), .C1(n4078), .C2(n6126), .A(n4658), 
        .ZN(n4645) );
  AOI22_X1 U2102 ( .A1(n6138), .A2(n4659), .B1(n6146), .B2(n4660), .ZN(n4658)
         );
  OAI221_X1 U2103 ( .B1(n4061), .B2(n6119), .C1(n4060), .C2(n6126), .A(n4624), 
        .ZN(n4611) );
  AOI22_X1 U2104 ( .A1(n6138), .A2(n4625), .B1(n6146), .B2(n4626), .ZN(n4624)
         );
  OAI221_X1 U2105 ( .B1(n4043), .B2(n6119), .C1(n4042), .C2(n6127), .A(n4590), 
        .ZN(n4577) );
  AOI22_X1 U2106 ( .A1(n6133), .A2(n4591), .B1(n6141), .B2(n4592), .ZN(n4590)
         );
  OAI221_X1 U2107 ( .B1(n4025), .B2(n6120), .C1(n4024), .C2(n6126), .A(n4556), 
        .ZN(n4543) );
  AOI22_X1 U2108 ( .A1(n6137), .A2(n4557), .B1(n6145), .B2(n4558), .ZN(n4556)
         );
  OAI221_X1 U2109 ( .B1(n4007), .B2(n6122), .C1(n4006), .C2(n6131), .A(n4522), 
        .ZN(n4509) );
  AOI22_X1 U2110 ( .A1(n6135), .A2(n4523), .B1(n6146), .B2(n4524), .ZN(n4522)
         );
  OAI221_X1 U2111 ( .B1(n3989), .B2(n6123), .C1(n3988), .C2(n6130), .A(n4488), 
        .ZN(n4475) );
  AOI22_X1 U2112 ( .A1(n6138), .A2(n4489), .B1(n6146), .B2(n4490), .ZN(n4488)
         );
  OAI221_X1 U2113 ( .B1(n3971), .B2(n6123), .C1(n3970), .C2(n6128), .A(n4454), 
        .ZN(n4441) );
  AOI22_X1 U2114 ( .A1(n6139), .A2(n4455), .B1(n6147), .B2(n4456), .ZN(n4454)
         );
  OAI221_X1 U2115 ( .B1(n3953), .B2(n6121), .C1(n3952), .C2(n6128), .A(n4420), 
        .ZN(n4407) );
  AOI22_X1 U2116 ( .A1(n6139), .A2(n4421), .B1(n6147), .B2(n4422), .ZN(n4420)
         );
  OAI221_X1 U2117 ( .B1(n3935), .B2(n6121), .C1(n3934), .C2(n6129), .A(n4386), 
        .ZN(n4373) );
  AOI22_X1 U2118 ( .A1(n6139), .A2(n4387), .B1(n6147), .B2(n4388), .ZN(n4386)
         );
  OAI221_X1 U2119 ( .B1(n3917), .B2(n6122), .C1(n3916), .C2(n6130), .A(n4352), 
        .ZN(n4339) );
  AOI22_X1 U2120 ( .A1(n6139), .A2(n4353), .B1(n6147), .B2(n4354), .ZN(n4352)
         );
  OAI221_X1 U2121 ( .B1(n3881), .B2(n6122), .C1(n3880), .C2(n6130), .A(n3708), 
        .ZN(n3695) );
  AOI22_X1 U2122 ( .A1(n6138), .A2(n3709), .B1(n6143), .B2(n3710), .ZN(n3708)
         );
  OAI221_X1 U2123 ( .B1(n3863), .B2(n6123), .C1(n3862), .C2(n6131), .A(n2649), 
        .ZN(n2636) );
  AOI22_X1 U2124 ( .A1(n6138), .A2(n2650), .B1(n6144), .B2(n2651), .ZN(n2649)
         );
  OAI221_X1 U2125 ( .B1(n2006), .B2(n6281), .C1(n65), .C2(n6289), .A(n4299), 
        .ZN(n3714) );
  AOI22_X1 U2126 ( .A1(n6293), .A2(n4300), .B1(n6302), .B2(n4301), .ZN(n4299)
         );
  OAI221_X1 U2127 ( .B1(n2306), .B2(n6153), .C1(n68), .C2(n6161), .A(n4315), 
        .ZN(n4306) );
  AOI22_X1 U2128 ( .A1(n6169), .A2(n4316), .B1(n6173), .B2(n4317), .ZN(n4315)
         );
  OAI221_X1 U2129 ( .B1(n2005), .B2(n6282), .C1(n44), .C2(n6291), .A(n2596), 
        .ZN(n2587) );
  AOI22_X1 U2130 ( .A1(n6294), .A2(n2597), .B1(n6301), .B2(n2598), .ZN(n2596)
         );
  OAI221_X1 U2131 ( .B1(n2305), .B2(n6154), .C1(n47), .C2(n6163), .A(n2612), 
        .ZN(n2603) );
  AOI22_X1 U2132 ( .A1(n6165), .A2(n2613), .B1(n6173), .B2(n2614), .ZN(n2612)
         );
  OAI221_X1 U2133 ( .B1(n2304), .B2(n6154), .C1(n40), .C2(n6162), .A(n2578), 
        .ZN(n2569) );
  AOI22_X1 U2134 ( .A1(n6165), .A2(n2579), .B1(n6174), .B2(n2580), .ZN(n2578)
         );
  OAI221_X1 U2135 ( .B1(n2000), .B2(n6282), .C1(n9), .C2(n6290), .A(n2426), 
        .ZN(n2417) );
  AOI22_X1 U2136 ( .A1(n6296), .A2(n2427), .B1(n6303), .B2(n2428), .ZN(n2426)
         );
  OAI221_X1 U2137 ( .B1(n2299), .B2(n6151), .C1(n5), .C2(n6160), .A(n2402), 
        .ZN(n2383) );
  AOI22_X1 U2138 ( .A1(n6168), .A2(n2404), .B1(n6177), .B2(n2406), .ZN(n2402)
         );
  OAI221_X1 U2139 ( .B1(n1984), .B2(n6280), .C1(n93), .C2(n6288), .A(n4435), 
        .ZN(n4426) );
  AOI22_X1 U2140 ( .A1(n6297), .A2(n4436), .B1(n6307), .B2(n4437), .ZN(n4435)
         );
  OAI221_X1 U2141 ( .B1(n2285), .B2(n6153), .C1(n96), .C2(n6160), .A(n4451), 
        .ZN(n4442) );
  AOI22_X1 U2142 ( .A1(n6171), .A2(n4452), .B1(n6179), .B2(n4453), .ZN(n4451)
         );
  OAI221_X1 U2143 ( .B1(n1983), .B2(n6281), .C1(n86), .C2(n6288), .A(n4401), 
        .ZN(n4392) );
  AOI22_X1 U2144 ( .A1(n6295), .A2(n4402), .B1(n6307), .B2(n4403), .ZN(n4401)
         );
  OAI221_X1 U2145 ( .B1(n2284), .B2(n6153), .C1(n89), .C2(n6160), .A(n4417), 
        .ZN(n4408) );
  AOI22_X1 U2146 ( .A1(n6171), .A2(n4418), .B1(n6179), .B2(n4419), .ZN(n4417)
         );
  OAI221_X1 U2147 ( .B1(n1982), .B2(n6281), .C1(n79), .C2(n6289), .A(n4367), 
        .ZN(n4358) );
  AOI22_X1 U2148 ( .A1(n6296), .A2(n4368), .B1(n6307), .B2(n4369), .ZN(n4367)
         );
  OAI221_X1 U2149 ( .B1(n2283), .B2(n6153), .C1(n82), .C2(n6161), .A(n4383), 
        .ZN(n4374) );
  AOI22_X1 U2150 ( .A1(n6171), .A2(n4384), .B1(n6179), .B2(n4385), .ZN(n4383)
         );
  OAI221_X1 U2151 ( .B1(n1981), .B2(n6283), .C1(n72), .C2(n6290), .A(n4333), 
        .ZN(n4324) );
  AOI22_X1 U2152 ( .A1(n6299), .A2(n4334), .B1(n6307), .B2(n4335), .ZN(n4333)
         );
  OAI221_X1 U2153 ( .B1(n2282), .B2(n6154), .C1(n75), .C2(n6162), .A(n4349), 
        .ZN(n4340) );
  AOI22_X1 U2154 ( .A1(n6171), .A2(n4350), .B1(n6179), .B2(n4351), .ZN(n4349)
         );
  OAI221_X1 U2155 ( .B1(n1980), .B2(n6283), .C1(n58), .C2(n6290), .A(n3689), 
        .ZN(n2655) );
  AOI22_X1 U2156 ( .A1(n6297), .A2(n3690), .B1(n6304), .B2(n3691), .ZN(n3689)
         );
  OAI221_X1 U2157 ( .B1(n2281), .B2(n6155), .C1(n61), .C2(n6162), .A(n3705), 
        .ZN(n3696) );
  AOI22_X1 U2158 ( .A1(n6165), .A2(n3706), .B1(n6176), .B2(n3707), .ZN(n3705)
         );
  OAI221_X1 U2159 ( .B1(n1979), .B2(n6282), .C1(n51), .C2(n6291), .A(n2630), 
        .ZN(n2621) );
  AOI22_X1 U2160 ( .A1(n6296), .A2(n2631), .B1(n6303), .B2(n2632), .ZN(n2630)
         );
  OAI221_X1 U2161 ( .B1(n2280), .B2(n6155), .C1(n54), .C2(n6163), .A(n2646), 
        .ZN(n2637) );
  AOI22_X1 U2162 ( .A1(n6166), .A2(n2647), .B1(n6175), .B2(n2648), .ZN(n2646)
         );
  OAI221_X1 U2163 ( .B1(n1937), .B2(n6249), .C1(n64), .C2(n6257), .A(n4302), 
        .ZN(n3713) );
  AOI22_X1 U2164 ( .A1(n6261), .A2(n4303), .B1(n6270), .B2(n4304), .ZN(n4302)
         );
  OAI221_X1 U2165 ( .B1(n1935), .B2(n6250), .C1(n43), .C2(n6259), .A(n2599), 
        .ZN(n2586) );
  AOI22_X1 U2166 ( .A1(n6262), .A2(n2600), .B1(n6269), .B2(n2601), .ZN(n2599)
         );
  OAI221_X1 U2167 ( .B1(n1925), .B2(n6251), .C1(n8), .C2(n6254), .A(n2429), 
        .ZN(n2416) );
  AOI22_X1 U2168 ( .A1(n6263), .A2(n2430), .B1(n6272), .B2(n2431), .ZN(n2429)
         );
  OAI221_X1 U2169 ( .B1(n1893), .B2(n6246), .C1(n99), .C2(n6258), .A(n4472), 
        .ZN(n4459) );
  AOI22_X1 U2170 ( .A1(n6267), .A2(n4473), .B1(n6274), .B2(n4474), .ZN(n4472)
         );
  OAI221_X1 U2171 ( .B1(n1891), .B2(n6248), .C1(n92), .C2(n6256), .A(n4438), 
        .ZN(n4425) );
  AOI22_X1 U2172 ( .A1(n6267), .A2(n4439), .B1(n6275), .B2(n4440), .ZN(n4438)
         );
  OAI221_X1 U2173 ( .B1(n1889), .B2(n6249), .C1(n85), .C2(n6256), .A(n4404), 
        .ZN(n4391) );
  AOI22_X1 U2174 ( .A1(n6267), .A2(n4405), .B1(n6275), .B2(n4406), .ZN(n4404)
         );
  OAI221_X1 U2175 ( .B1(n1887), .B2(n6249), .C1(n78), .C2(n6257), .A(n4370), 
        .ZN(n4357) );
  AOI22_X1 U2176 ( .A1(n6267), .A2(n4371), .B1(n6275), .B2(n4372), .ZN(n4370)
         );
  OAI221_X1 U2177 ( .B1(n1885), .B2(n6251), .C1(n71), .C2(n6258), .A(n4336), 
        .ZN(n4323) );
  AOI22_X1 U2178 ( .A1(n6267), .A2(n4337), .B1(n6275), .B2(n4338), .ZN(n4336)
         );
  OAI221_X1 U2179 ( .B1(n1883), .B2(n6251), .C1(n57), .C2(n6258), .A(n3692), 
        .ZN(n2654) );
  AOI22_X1 U2180 ( .A1(n6264), .A2(n3693), .B1(n6271), .B2(n3694), .ZN(n3692)
         );
  OAI221_X1 U2181 ( .B1(n1881), .B2(n6250), .C1(n50), .C2(n6259), .A(n2633), 
        .ZN(n2620) );
  AOI22_X1 U2182 ( .A1(n6263), .A2(n2634), .B1(n6271), .B2(n2635), .ZN(n2633)
         );
  NOR3_X1 U2183 ( .A1(n5726), .A2(n5082), .A3(n5727), .ZN(n5725) );
  XNOR2_X1 U2184 ( .A(n2340), .B(ADD_RD2[1]), .ZN(n5726) );
  XNOR2_X1 U2185 ( .A(ADD_WR[4]), .B(n5075), .ZN(n5727) );
  AOI211_X1 U2186 ( .C1(n5713), .C2(n5714), .A(n6736), .B(n2158), .ZN(N4192)
         );
  NAND4_X1 U2187 ( .A1(n5716), .A2(n5717), .A3(n5718), .A4(n5719), .ZN(n5714)
         );
  NAND4_X1 U2188 ( .A1(n5722), .A2(n5723), .A3(n5724), .A4(n5725), .ZN(n5713)
         );
  XNOR2_X1 U2189 ( .A(ADD_RD1[2]), .B(ADD_WR[2]), .ZN(n5716) );
  INV_X1 U2190 ( .A(ADD_RD2[4]), .ZN(n5075) );
  NOR2_X1 U2191 ( .A1(n2158), .A2(ADD_WR[4]), .ZN(n1976) );
  OAI22_X1 U2192 ( .A1(n6356), .A2(n6629), .B1(net86667), .B2(n6348), .ZN(
        n2657) );
  OAI22_X1 U2193 ( .A1(n6364), .A2(n6703), .B1(net86723), .B2(n2345), .ZN(
        n2713) );
  OAI22_X1 U2194 ( .A1(n6365), .A2(n6706), .B1(net86724), .B2(n6359), .ZN(
        n2714) );
  OAI22_X1 U2195 ( .A1(n6365), .A2(n6709), .B1(net86725), .B2(n6359), .ZN(
        n2715) );
  OAI22_X1 U2196 ( .A1(n6365), .A2(n6712), .B1(net86726), .B2(n6359), .ZN(
        n2716) );
  OAI22_X1 U2197 ( .A1(n6365), .A2(n6715), .B1(net86727), .B2(n6359), .ZN(
        n2717) );
  OAI22_X1 U2198 ( .A1(n6365), .A2(n6718), .B1(net86728), .B2(n2345), .ZN(
        n2718) );
  OAI22_X1 U2199 ( .A1(n6366), .A2(n6721), .B1(net86729), .B2(n6359), .ZN(
        n2719) );
  OAI22_X1 U2200 ( .A1(n6366), .A2(n6733), .B1(net86730), .B2(n2345), .ZN(
        n2720) );
  OAI22_X1 U2201 ( .A1(n6373), .A2(n6703), .B1(n4007), .B2(n2343), .ZN(n2745)
         );
  OAI22_X1 U2202 ( .A1(n6374), .A2(n6706), .B1(n3989), .B2(n6368), .ZN(n2746)
         );
  OAI22_X1 U2203 ( .A1(n6374), .A2(n6709), .B1(n3971), .B2(n6368), .ZN(n2747)
         );
  OAI22_X1 U2204 ( .A1(n6374), .A2(n6712), .B1(n3953), .B2(n6368), .ZN(n2748)
         );
  OAI22_X1 U2205 ( .A1(n6374), .A2(n6715), .B1(n3935), .B2(n6368), .ZN(n2749)
         );
  OAI22_X1 U2206 ( .A1(n6374), .A2(n6718), .B1(n3917), .B2(n2343), .ZN(n2750)
         );
  OAI22_X1 U2207 ( .A1(n6375), .A2(n6721), .B1(n3881), .B2(n6368), .ZN(n2751)
         );
  OAI22_X1 U2208 ( .A1(n6375), .A2(n6733), .B1(n3863), .B2(n2343), .ZN(n2752)
         );
  OAI22_X1 U2209 ( .A1(n6382), .A2(n6703), .B1(n4006), .B2(n2338), .ZN(n2777)
         );
  OAI22_X1 U2210 ( .A1(n6383), .A2(n6706), .B1(n3988), .B2(n6377), .ZN(n2778)
         );
  OAI22_X1 U2211 ( .A1(n6383), .A2(n6709), .B1(n3970), .B2(n6377), .ZN(n2779)
         );
  OAI22_X1 U2212 ( .A1(n6383), .A2(n6712), .B1(n3952), .B2(n6377), .ZN(n2780)
         );
  OAI22_X1 U2213 ( .A1(n6383), .A2(n6715), .B1(n3934), .B2(n6377), .ZN(n2781)
         );
  OAI22_X1 U2214 ( .A1(n6383), .A2(n6718), .B1(n3916), .B2(n2338), .ZN(n2782)
         );
  OAI22_X1 U2215 ( .A1(n6384), .A2(n6721), .B1(n3880), .B2(n6377), .ZN(n2783)
         );
  OAI22_X1 U2216 ( .A1(n6384), .A2(n6733), .B1(n3862), .B2(n2338), .ZN(n2784)
         );
  OAI22_X1 U2217 ( .A1(n6391), .A2(n6703), .B1(net86755), .B2(n2336), .ZN(
        n2809) );
  OAI22_X1 U2218 ( .A1(n6392), .A2(n6706), .B1(net86756), .B2(n6386), .ZN(
        n2810) );
  OAI22_X1 U2219 ( .A1(n6392), .A2(n6709), .B1(net86757), .B2(n6386), .ZN(
        n2811) );
  OAI22_X1 U2220 ( .A1(n6392), .A2(n6712), .B1(net86758), .B2(n6386), .ZN(
        n2812) );
  OAI22_X1 U2221 ( .A1(n6392), .A2(n6715), .B1(net86759), .B2(n6386), .ZN(
        n2813) );
  OAI22_X1 U2222 ( .A1(n6392), .A2(n6718), .B1(net86760), .B2(n2336), .ZN(
        n2814) );
  OAI22_X1 U2223 ( .A1(n6393), .A2(n6721), .B1(net86761), .B2(n6386), .ZN(
        n2815) );
  OAI22_X1 U2224 ( .A1(n6393), .A2(n6733), .B1(net86762), .B2(n2336), .ZN(
        n2816) );
  OAI22_X1 U2225 ( .A1(n6400), .A2(n6703), .B1(net86787), .B2(n2334), .ZN(
        n2841) );
  OAI22_X1 U2226 ( .A1(n6401), .A2(n6706), .B1(net86788), .B2(n6395), .ZN(
        n2842) );
  OAI22_X1 U2227 ( .A1(n6401), .A2(n6709), .B1(net86789), .B2(n6395), .ZN(
        n2843) );
  OAI22_X1 U2228 ( .A1(n6401), .A2(n6712), .B1(net86790), .B2(n6395), .ZN(
        n2844) );
  OAI22_X1 U2229 ( .A1(n6401), .A2(n6715), .B1(net86791), .B2(n6395), .ZN(
        n2845) );
  OAI22_X1 U2230 ( .A1(n6401), .A2(n6718), .B1(net86792), .B2(n2334), .ZN(
        n2846) );
  OAI22_X1 U2231 ( .A1(n6402), .A2(n6721), .B1(net86793), .B2(n6395), .ZN(
        n2847) );
  OAI22_X1 U2232 ( .A1(n6402), .A2(n6733), .B1(net86794), .B2(n2334), .ZN(
        n2848) );
  OAI22_X1 U2233 ( .A1(n6427), .A2(n6702), .B1(net86819), .B2(n2277), .ZN(
        n2937) );
  OAI22_X1 U2234 ( .A1(n6428), .A2(n6705), .B1(net86820), .B2(n6422), .ZN(
        n2938) );
  OAI22_X1 U2235 ( .A1(n6428), .A2(n6708), .B1(net86821), .B2(n6422), .ZN(
        n2939) );
  OAI22_X1 U2236 ( .A1(n6428), .A2(n6711), .B1(net86822), .B2(n6422), .ZN(
        n2940) );
  OAI22_X1 U2237 ( .A1(n6428), .A2(n6714), .B1(net86823), .B2(n6422), .ZN(
        n2941) );
  OAI22_X1 U2238 ( .A1(n6428), .A2(n6717), .B1(net86824), .B2(n2277), .ZN(
        n2942) );
  OAI22_X1 U2239 ( .A1(n6429), .A2(n6720), .B1(net86825), .B2(n6422), .ZN(
        n2943) );
  OAI22_X1 U2240 ( .A1(n6429), .A2(n6732), .B1(net86826), .B2(n2277), .ZN(
        n2944) );
  OAI22_X1 U2241 ( .A1(n6436), .A2(n6702), .B1(net86851), .B2(n2275), .ZN(
        n2969) );
  OAI22_X1 U2242 ( .A1(n6437), .A2(n6705), .B1(net86852), .B2(n6431), .ZN(
        n2970) );
  OAI22_X1 U2243 ( .A1(n6437), .A2(n6708), .B1(net86853), .B2(n6431), .ZN(
        n2971) );
  OAI22_X1 U2244 ( .A1(n6437), .A2(n6711), .B1(net86854), .B2(n6431), .ZN(
        n2972) );
  OAI22_X1 U2245 ( .A1(n6437), .A2(n6714), .B1(net86855), .B2(n6431), .ZN(
        n2973) );
  OAI22_X1 U2246 ( .A1(n6437), .A2(n6717), .B1(net86856), .B2(n2275), .ZN(
        n2974) );
  OAI22_X1 U2247 ( .A1(n6438), .A2(n6720), .B1(net86857), .B2(n6431), .ZN(
        n2975) );
  OAI22_X1 U2248 ( .A1(n6438), .A2(n6732), .B1(net86858), .B2(n2275), .ZN(
        n2976) );
  OAI22_X1 U2249 ( .A1(n6463), .A2(n6702), .B1(net86883), .B2(n2217), .ZN(
        n3065) );
  OAI22_X1 U2250 ( .A1(n6464), .A2(n6705), .B1(net86884), .B2(n6458), .ZN(
        n3066) );
  OAI22_X1 U2251 ( .A1(n6464), .A2(n6708), .B1(net86885), .B2(n6458), .ZN(
        n3067) );
  OAI22_X1 U2252 ( .A1(n6464), .A2(n6711), .B1(net86886), .B2(n6458), .ZN(
        n3068) );
  OAI22_X1 U2253 ( .A1(n6464), .A2(n6714), .B1(net86887), .B2(n6458), .ZN(
        n3069) );
  OAI22_X1 U2254 ( .A1(n6464), .A2(n6717), .B1(net86888), .B2(n2217), .ZN(
        n3070) );
  OAI22_X1 U2255 ( .A1(n6465), .A2(n6720), .B1(net86889), .B2(n6458), .ZN(
        n3071) );
  OAI22_X1 U2256 ( .A1(n6465), .A2(n6732), .B1(net86890), .B2(n2217), .ZN(
        n3072) );
  OAI22_X1 U2257 ( .A1(n6472), .A2(n6702), .B1(net86915), .B2(n2215), .ZN(
        n3097) );
  OAI22_X1 U2258 ( .A1(n6473), .A2(n6705), .B1(net86916), .B2(n6467), .ZN(
        n3098) );
  OAI22_X1 U2259 ( .A1(n6473), .A2(n6708), .B1(net86917), .B2(n6467), .ZN(
        n3099) );
  OAI22_X1 U2260 ( .A1(n6473), .A2(n6711), .B1(net86918), .B2(n6467), .ZN(
        n3100) );
  OAI22_X1 U2261 ( .A1(n6473), .A2(n6714), .B1(net86919), .B2(n6467), .ZN(
        n3101) );
  OAI22_X1 U2262 ( .A1(n6473), .A2(n6717), .B1(net86920), .B2(n2215), .ZN(
        n3102) );
  OAI22_X1 U2263 ( .A1(n6474), .A2(n6720), .B1(net86921), .B2(n6467), .ZN(
        n3103) );
  OAI22_X1 U2264 ( .A1(n6474), .A2(n6732), .B1(net86922), .B2(n2215), .ZN(
        n3104) );
  OAI22_X1 U2265 ( .A1(n6499), .A2(n6702), .B1(net86947), .B2(n2157), .ZN(
        n3193) );
  OAI22_X1 U2266 ( .A1(n6500), .A2(n6705), .B1(net86948), .B2(n6494), .ZN(
        n3194) );
  OAI22_X1 U2267 ( .A1(n6500), .A2(n6708), .B1(net86949), .B2(n6494), .ZN(
        n3195) );
  OAI22_X1 U2268 ( .A1(n6500), .A2(n6711), .B1(net86950), .B2(n6494), .ZN(
        n3196) );
  OAI22_X1 U2269 ( .A1(n6500), .A2(n6714), .B1(net86951), .B2(n6494), .ZN(
        n3197) );
  OAI22_X1 U2270 ( .A1(n6500), .A2(n6717), .B1(net86952), .B2(n2157), .ZN(
        n3198) );
  OAI22_X1 U2271 ( .A1(n6501), .A2(n6720), .B1(net86953), .B2(n6494), .ZN(
        n3199) );
  OAI22_X1 U2272 ( .A1(n6501), .A2(n6732), .B1(net86954), .B2(n2157), .ZN(
        n3200) );
  OAI22_X1 U2273 ( .A1(n6508), .A2(n6702), .B1(net86979), .B2(n2155), .ZN(
        n3225) );
  OAI22_X1 U2274 ( .A1(n6509), .A2(n6705), .B1(net86980), .B2(n6503), .ZN(
        n3226) );
  OAI22_X1 U2275 ( .A1(n6509), .A2(n6708), .B1(net86981), .B2(n6503), .ZN(
        n3227) );
  OAI22_X1 U2276 ( .A1(n6509), .A2(n6711), .B1(net86982), .B2(n6503), .ZN(
        n3228) );
  OAI22_X1 U2277 ( .A1(n6509), .A2(n6714), .B1(net86983), .B2(n6503), .ZN(
        n3229) );
  OAI22_X1 U2278 ( .A1(n6509), .A2(n6717), .B1(net86984), .B2(n2155), .ZN(
        n3230) );
  OAI22_X1 U2279 ( .A1(n6510), .A2(n6720), .B1(net86985), .B2(n6503), .ZN(
        n3231) );
  OAI22_X1 U2280 ( .A1(n6510), .A2(n6732), .B1(net86986), .B2(n2155), .ZN(
        n3232) );
  OAI22_X1 U2281 ( .A1(n6535), .A2(n6701), .B1(net87011), .B2(n2098), .ZN(
        n3321) );
  OAI22_X1 U2282 ( .A1(n6536), .A2(n6704), .B1(net87012), .B2(n6530), .ZN(
        n3322) );
  OAI22_X1 U2283 ( .A1(n6536), .A2(n6707), .B1(net87013), .B2(n6530), .ZN(
        n3323) );
  OAI22_X1 U2284 ( .A1(n6536), .A2(n6710), .B1(net87014), .B2(n6530), .ZN(
        n3324) );
  OAI22_X1 U2285 ( .A1(n6536), .A2(n6713), .B1(net87015), .B2(n6530), .ZN(
        n3325) );
  OAI22_X1 U2286 ( .A1(n6536), .A2(n6716), .B1(net87016), .B2(n2098), .ZN(
        n3326) );
  OAI22_X1 U2287 ( .A1(n6537), .A2(n6719), .B1(net87017), .B2(n6530), .ZN(
        n3327) );
  OAI22_X1 U2288 ( .A1(n6537), .A2(n6731), .B1(net87018), .B2(n2098), .ZN(
        n3328) );
  OAI22_X1 U2289 ( .A1(n6544), .A2(n6701), .B1(net87043), .B2(n2096), .ZN(
        n3353) );
  OAI22_X1 U2290 ( .A1(n6545), .A2(n6704), .B1(net87044), .B2(n6539), .ZN(
        n3354) );
  OAI22_X1 U2291 ( .A1(n6545), .A2(n6707), .B1(net87045), .B2(n6539), .ZN(
        n3355) );
  OAI22_X1 U2292 ( .A1(n6545), .A2(n6710), .B1(net87046), .B2(n6539), .ZN(
        n3356) );
  OAI22_X1 U2293 ( .A1(n6545), .A2(n6713), .B1(net87047), .B2(n6539), .ZN(
        n3357) );
  OAI22_X1 U2294 ( .A1(n6545), .A2(n6716), .B1(net87048), .B2(n2096), .ZN(
        n3358) );
  OAI22_X1 U2295 ( .A1(n6546), .A2(n6719), .B1(net87049), .B2(n6539), .ZN(
        n3359) );
  OAI22_X1 U2296 ( .A1(n6546), .A2(n6731), .B1(net87050), .B2(n2096), .ZN(
        n3360) );
  OAI22_X1 U2297 ( .A1(n6571), .A2(n6701), .B1(net87075), .B2(n2037), .ZN(
        n3449) );
  OAI22_X1 U2298 ( .A1(n6572), .A2(n6704), .B1(net87076), .B2(n6566), .ZN(
        n3450) );
  OAI22_X1 U2299 ( .A1(n6572), .A2(n6707), .B1(net87077), .B2(n6566), .ZN(
        n3451) );
  OAI22_X1 U2300 ( .A1(n6572), .A2(n6710), .B1(net87078), .B2(n6566), .ZN(
        n3452) );
  OAI22_X1 U2301 ( .A1(n6572), .A2(n6713), .B1(net87079), .B2(n6566), .ZN(
        n3453) );
  OAI22_X1 U2302 ( .A1(n6572), .A2(n6716), .B1(net87080), .B2(n2037), .ZN(
        n3454) );
  OAI22_X1 U2303 ( .A1(n6573), .A2(n6719), .B1(net87081), .B2(n6566), .ZN(
        n3455) );
  OAI22_X1 U2304 ( .A1(n6573), .A2(n6731), .B1(net87082), .B2(n2037), .ZN(
        n3456) );
  OAI22_X1 U2305 ( .A1(n6580), .A2(n6701), .B1(net87107), .B2(n2035), .ZN(
        n3481) );
  OAI22_X1 U2306 ( .A1(n6581), .A2(n6704), .B1(net87108), .B2(n6575), .ZN(
        n3482) );
  OAI22_X1 U2307 ( .A1(n6581), .A2(n6707), .B1(net87109), .B2(n6575), .ZN(
        n3483) );
  OAI22_X1 U2308 ( .A1(n6581), .A2(n6710), .B1(net87110), .B2(n6575), .ZN(
        n3484) );
  OAI22_X1 U2309 ( .A1(n6581), .A2(n6713), .B1(net87111), .B2(n6575), .ZN(
        n3485) );
  OAI22_X1 U2310 ( .A1(n6581), .A2(n6716), .B1(net87112), .B2(n2035), .ZN(
        n3486) );
  OAI22_X1 U2311 ( .A1(n6582), .A2(n6719), .B1(net87113), .B2(n6575), .ZN(
        n3487) );
  OAI22_X1 U2312 ( .A1(n6582), .A2(n6731), .B1(net87114), .B2(n2035), .ZN(
        n3488) );
  OAI22_X1 U2313 ( .A1(n6607), .A2(n6701), .B1(net87139), .B2(n1972), .ZN(
        n3577) );
  OAI22_X1 U2314 ( .A1(n6608), .A2(n6704), .B1(net87140), .B2(n6602), .ZN(
        n3578) );
  OAI22_X1 U2315 ( .A1(n6608), .A2(n6707), .B1(net87141), .B2(n6602), .ZN(
        n3579) );
  OAI22_X1 U2316 ( .A1(n6608), .A2(n6710), .B1(net87142), .B2(n6602), .ZN(
        n3580) );
  OAI22_X1 U2317 ( .A1(n6608), .A2(n6713), .B1(net87143), .B2(n6602), .ZN(
        n3581) );
  OAI22_X1 U2318 ( .A1(n6608), .A2(n6716), .B1(net87144), .B2(n1972), .ZN(
        n3582) );
  OAI22_X1 U2319 ( .A1(n6609), .A2(n6719), .B1(net87145), .B2(n6602), .ZN(
        n3583) );
  OAI22_X1 U2320 ( .A1(n6609), .A2(n6731), .B1(net87146), .B2(n1972), .ZN(
        n3584) );
  OAI22_X1 U2321 ( .A1(n6616), .A2(n6701), .B1(net87171), .B2(n1969), .ZN(
        n3609) );
  OAI22_X1 U2322 ( .A1(n6617), .A2(n6704), .B1(net87172), .B2(n6611), .ZN(
        n3610) );
  OAI22_X1 U2323 ( .A1(n6617), .A2(n6707), .B1(net87173), .B2(n6611), .ZN(
        n3611) );
  OAI22_X1 U2324 ( .A1(n6617), .A2(n6710), .B1(net87174), .B2(n6611), .ZN(
        n3612) );
  OAI22_X1 U2325 ( .A1(n6617), .A2(n6713), .B1(net87175), .B2(n6611), .ZN(
        n3613) );
  OAI22_X1 U2326 ( .A1(n6617), .A2(n6716), .B1(net87176), .B2(n1969), .ZN(
        n3614) );
  OAI22_X1 U2327 ( .A1(n6618), .A2(n6719), .B1(net87177), .B2(n6611), .ZN(
        n3615) );
  OAI22_X1 U2328 ( .A1(n6618), .A2(n6731), .B1(net87178), .B2(n1969), .ZN(
        n3616) );
  OAI22_X1 U2329 ( .A1(net86687), .A2(n6348), .B1(n6351), .B2(n6691), .ZN(
        n2677) );
  OAI22_X1 U2330 ( .A1(net86688), .A2(n6348), .B1(n6351), .B2(n6694), .ZN(
        n2678) );
  OAI22_X1 U2331 ( .A1(net86689), .A2(n6348), .B1(n6351), .B2(n6697), .ZN(
        n2679) );
  OAI22_X1 U2332 ( .A1(net86690), .A2(n6348), .B1(n6351), .B2(n6700), .ZN(
        n2680) );
  OAI22_X1 U2333 ( .A1(net86691), .A2(n6348), .B1(n6350), .B2(n6703), .ZN(
        n2681) );
  OAI22_X1 U2334 ( .A1(net86692), .A2(n6348), .B1(n6350), .B2(n6706), .ZN(
        n2682) );
  OAI22_X1 U2335 ( .A1(net86693), .A2(n6348), .B1(n6350), .B2(n6709), .ZN(
        n2683) );
  OAI22_X1 U2336 ( .A1(net86694), .A2(n6348), .B1(n6350), .B2(n6712), .ZN(
        n2684) );
  OAI22_X1 U2337 ( .A1(net86695), .A2(n6348), .B1(n6349), .B2(n6715), .ZN(
        n2685) );
  OAI22_X1 U2338 ( .A1(net86696), .A2(n6348), .B1(n6349), .B2(n6718), .ZN(
        n2686) );
  OAI22_X1 U2339 ( .A1(net86697), .A2(n6348), .B1(n6349), .B2(n6721), .ZN(
        n2687) );
  OAI22_X1 U2340 ( .A1(net86698), .A2(n6348), .B1(n6349), .B2(n6733), .ZN(
        n2688) );
  OAI22_X1 U2341 ( .A1(net86668), .A2(n2346), .B1(n6356), .B2(n6634), .ZN(
        n2658) );
  OAI22_X1 U2342 ( .A1(net86669), .A2(n6348), .B1(n6356), .B2(n6637), .ZN(
        n2659) );
  OAI22_X1 U2343 ( .A1(net86670), .A2(n6348), .B1(n6356), .B2(n6640), .ZN(
        n2660) );
  OAI22_X1 U2344 ( .A1(net86671), .A2(n6348), .B1(n6355), .B2(n6643), .ZN(
        n2661) );
  OAI22_X1 U2345 ( .A1(net86672), .A2(n2346), .B1(n6355), .B2(n6646), .ZN(
        n2662) );
  OAI22_X1 U2346 ( .A1(net86673), .A2(n2346), .B1(n6355), .B2(n6649), .ZN(
        n2663) );
  OAI22_X1 U2347 ( .A1(net86674), .A2(n2346), .B1(n6355), .B2(n6652), .ZN(
        n2664) );
  OAI22_X1 U2348 ( .A1(net86675), .A2(n6348), .B1(n6354), .B2(n6655), .ZN(
        n2665) );
  OAI22_X1 U2349 ( .A1(net86676), .A2(n6348), .B1(n6354), .B2(n6658), .ZN(
        n2666) );
  OAI22_X1 U2350 ( .A1(net86677), .A2(n2346), .B1(n6354), .B2(n6661), .ZN(
        n2667) );
  OAI22_X1 U2351 ( .A1(net86678), .A2(n6348), .B1(n6354), .B2(n6664), .ZN(
        n2668) );
  OAI22_X1 U2352 ( .A1(net86679), .A2(n2346), .B1(n6353), .B2(n6667), .ZN(
        n2669) );
  OAI22_X1 U2353 ( .A1(net86680), .A2(n2346), .B1(n6353), .B2(n6670), .ZN(
        n2670) );
  OAI22_X1 U2354 ( .A1(net86681), .A2(n2346), .B1(n6353), .B2(n6673), .ZN(
        n2671) );
  OAI22_X1 U2355 ( .A1(net86682), .A2(n6348), .B1(n6353), .B2(n6676), .ZN(
        n2672) );
  OAI22_X1 U2356 ( .A1(net86683), .A2(n2346), .B1(n6352), .B2(n6679), .ZN(
        n2673) );
  OAI22_X1 U2357 ( .A1(net86684), .A2(n2346), .B1(n6352), .B2(n6682), .ZN(
        n2674) );
  OAI22_X1 U2358 ( .A1(net86685), .A2(n2346), .B1(n6352), .B2(n6685), .ZN(
        n2675) );
  OAI22_X1 U2359 ( .A1(net86686), .A2(n6348), .B1(n6352), .B2(n6688), .ZN(
        n2676) );
  OAI22_X1 U2360 ( .A1(n6369), .A2(n6629), .B1(n4295), .B2(n6368), .ZN(n2721)
         );
  OAI22_X1 U2361 ( .A1(n6369), .A2(n6634), .B1(n4097), .B2(n6368), .ZN(n2722)
         );
  OAI22_X1 U2362 ( .A1(n6369), .A2(n6637), .B1(n3899), .B2(n6368), .ZN(n2723)
         );
  OAI22_X1 U2363 ( .A1(n6369), .A2(n6640), .B1(n3845), .B2(n6368), .ZN(n2724)
         );
  OAI22_X1 U2364 ( .A1(n6369), .A2(n6643), .B1(n3827), .B2(n6368), .ZN(n2725)
         );
  OAI22_X1 U2365 ( .A1(n6370), .A2(n6646), .B1(n3809), .B2(n6368), .ZN(n2726)
         );
  OAI22_X1 U2366 ( .A1(n6370), .A2(n6649), .B1(n3791), .B2(n6368), .ZN(n2727)
         );
  OAI22_X1 U2367 ( .A1(n6370), .A2(n6652), .B1(n3773), .B2(n6368), .ZN(n2728)
         );
  OAI22_X1 U2368 ( .A1(n6370), .A2(n6655), .B1(n3755), .B2(n6368), .ZN(n2729)
         );
  OAI22_X1 U2369 ( .A1(n6370), .A2(n6658), .B1(n3737), .B2(n6368), .ZN(n2730)
         );
  OAI22_X1 U2370 ( .A1(n6371), .A2(n6661), .B1(n4277), .B2(n6368), .ZN(n2731)
         );
  OAI22_X1 U2371 ( .A1(n6371), .A2(n6664), .B1(n4259), .B2(n6368), .ZN(n2732)
         );
  OAI22_X1 U2372 ( .A1(n6371), .A2(n6667), .B1(n4241), .B2(n2343), .ZN(n2733)
         );
  OAI22_X1 U2373 ( .A1(n6371), .A2(n6670), .B1(n4223), .B2(n2343), .ZN(n2734)
         );
  OAI22_X1 U2374 ( .A1(n6371), .A2(n6673), .B1(n4205), .B2(n2343), .ZN(n2735)
         );
  OAI22_X1 U2375 ( .A1(n6372), .A2(n6676), .B1(n4187), .B2(n2343), .ZN(n2736)
         );
  OAI22_X1 U2376 ( .A1(n6372), .A2(n6679), .B1(n4169), .B2(n2343), .ZN(n2737)
         );
  OAI22_X1 U2377 ( .A1(n6372), .A2(n6682), .B1(n4151), .B2(n2343), .ZN(n2738)
         );
  OAI22_X1 U2378 ( .A1(n6372), .A2(n6685), .B1(n4133), .B2(n2343), .ZN(n2739)
         );
  OAI22_X1 U2379 ( .A1(n6372), .A2(n6688), .B1(n4115), .B2(n2343), .ZN(n2740)
         );
  OAI22_X1 U2380 ( .A1(n6373), .A2(n6691), .B1(n4079), .B2(n6368), .ZN(n2741)
         );
  OAI22_X1 U2381 ( .A1(n6373), .A2(n6694), .B1(n4061), .B2(n6368), .ZN(n2742)
         );
  OAI22_X1 U2382 ( .A1(n6373), .A2(n6697), .B1(n4043), .B2(n6368), .ZN(n2743)
         );
  OAI22_X1 U2383 ( .A1(n6373), .A2(n6700), .B1(n4025), .B2(n6368), .ZN(n2744)
         );
  OAI22_X1 U2384 ( .A1(n6414), .A2(n6629), .B1(n446), .B2(n6413), .ZN(n2881)
         );
  OAI22_X1 U2385 ( .A1(n6416), .A2(n6661), .B1(n439), .B2(n6413), .ZN(n2891)
         );
  OAI22_X1 U2386 ( .A1(n6416), .A2(n6664), .B1(n432), .B2(n6413), .ZN(n2892)
         );
  OAI22_X1 U2387 ( .A1(n6416), .A2(n6667), .B1(n425), .B2(n6413), .ZN(n2893)
         );
  OAI22_X1 U2388 ( .A1(n6441), .A2(n6629), .B1(n448), .B2(n6440), .ZN(n2977)
         );
  OAI22_X1 U2389 ( .A1(n6443), .A2(n6660), .B1(n441), .B2(n6440), .ZN(n2987)
         );
  OAI22_X1 U2390 ( .A1(n6443), .A2(n6663), .B1(n434), .B2(n6440), .ZN(n2988)
         );
  OAI22_X1 U2391 ( .A1(n6443), .A2(n6666), .B1(n427), .B2(n6440), .ZN(n2989)
         );
  OAI22_X1 U2392 ( .A1(n6477), .A2(n6630), .B1(n447), .B2(n6476), .ZN(n3105)
         );
  OAI22_X1 U2393 ( .A1(n6479), .A2(n6660), .B1(n440), .B2(n6476), .ZN(n3115)
         );
  OAI22_X1 U2394 ( .A1(n6479), .A2(n6663), .B1(n433), .B2(n6476), .ZN(n3116)
         );
  OAI22_X1 U2395 ( .A1(n6479), .A2(n6666), .B1(n426), .B2(n6476), .ZN(n3117)
         );
  OAI22_X1 U2396 ( .A1(n6522), .A2(n6630), .B1(n445), .B2(n6521), .ZN(n3265)
         );
  OAI22_X1 U2397 ( .A1(n6524), .A2(n6660), .B1(n438), .B2(n6521), .ZN(n3275)
         );
  OAI22_X1 U2398 ( .A1(n6524), .A2(n6663), .B1(n431), .B2(n6521), .ZN(n3276)
         );
  OAI22_X1 U2399 ( .A1(n6524), .A2(n6666), .B1(n424), .B2(n6521), .ZN(n3277)
         );
  OAI22_X1 U2400 ( .A1(n6558), .A2(n6630), .B1(n444), .B2(n6557), .ZN(n3393)
         );
  OAI22_X1 U2401 ( .A1(n6560), .A2(n6659), .B1(n437), .B2(n6557), .ZN(n3403)
         );
  OAI22_X1 U2402 ( .A1(n6560), .A2(n6662), .B1(n430), .B2(n6557), .ZN(n3404)
         );
  OAI22_X1 U2403 ( .A1(n6560), .A2(n6665), .B1(n423), .B2(n6557), .ZN(n3405)
         );
  OAI22_X1 U2404 ( .A1(n6594), .A2(n6631), .B1(n443), .B2(n6593), .ZN(n3521)
         );
  OAI22_X1 U2405 ( .A1(n6596), .A2(n6659), .B1(n436), .B2(n6593), .ZN(n3531)
         );
  OAI22_X1 U2406 ( .A1(n6596), .A2(n6662), .B1(n429), .B2(n6593), .ZN(n3532)
         );
  OAI22_X1 U2407 ( .A1(n6723), .A2(n6631), .B1(n442), .B2(n6722), .ZN(n3649)
         );
  OAI22_X1 U2408 ( .A1(n6725), .A2(n6659), .B1(n435), .B2(n6722), .ZN(n3659)
         );
  OAI22_X1 U2409 ( .A1(n6725), .A2(n6662), .B1(n428), .B2(n6722), .ZN(n3660)
         );
  OAI22_X1 U2410 ( .A1(n6360), .A2(n6629), .B1(net86699), .B2(n6359), .ZN(
        n2689) );
  OAI22_X1 U2411 ( .A1(n6360), .A2(n6634), .B1(net86700), .B2(n6359), .ZN(
        n2690) );
  OAI22_X1 U2412 ( .A1(n6360), .A2(n6637), .B1(net86701), .B2(n6359), .ZN(
        n2691) );
  OAI22_X1 U2413 ( .A1(n6360), .A2(n6640), .B1(net86702), .B2(n6359), .ZN(
        n2692) );
  OAI22_X1 U2414 ( .A1(n6360), .A2(n6643), .B1(net86703), .B2(n6359), .ZN(
        n2693) );
  OAI22_X1 U2415 ( .A1(n6361), .A2(n6646), .B1(net86704), .B2(n6359), .ZN(
        n2694) );
  OAI22_X1 U2416 ( .A1(n6361), .A2(n6649), .B1(net86705), .B2(n6359), .ZN(
        n2695) );
  OAI22_X1 U2417 ( .A1(n6361), .A2(n6652), .B1(net86706), .B2(n6359), .ZN(
        n2696) );
  OAI22_X1 U2418 ( .A1(n6361), .A2(n6655), .B1(net86707), .B2(n6359), .ZN(
        n2697) );
  OAI22_X1 U2419 ( .A1(n6361), .A2(n6658), .B1(net86708), .B2(n6359), .ZN(
        n2698) );
  OAI22_X1 U2420 ( .A1(n6362), .A2(n6661), .B1(net86709), .B2(n6359), .ZN(
        n2699) );
  OAI22_X1 U2421 ( .A1(n6362), .A2(n6664), .B1(net86710), .B2(n6359), .ZN(
        n2700) );
  OAI22_X1 U2422 ( .A1(n6362), .A2(n6667), .B1(net86711), .B2(n2345), .ZN(
        n2701) );
  OAI22_X1 U2423 ( .A1(n6362), .A2(n6670), .B1(net86712), .B2(n2345), .ZN(
        n2702) );
  OAI22_X1 U2424 ( .A1(n6362), .A2(n6673), .B1(net86713), .B2(n2345), .ZN(
        n2703) );
  OAI22_X1 U2425 ( .A1(n6363), .A2(n6676), .B1(net86714), .B2(n2345), .ZN(
        n2704) );
  OAI22_X1 U2426 ( .A1(n6363), .A2(n6679), .B1(net86715), .B2(n2345), .ZN(
        n2705) );
  OAI22_X1 U2427 ( .A1(n6363), .A2(n6682), .B1(net86716), .B2(n2345), .ZN(
        n2706) );
  OAI22_X1 U2428 ( .A1(n6363), .A2(n6685), .B1(net86717), .B2(n2345), .ZN(
        n2707) );
  OAI22_X1 U2429 ( .A1(n6363), .A2(n6688), .B1(net86718), .B2(n2345), .ZN(
        n2708) );
  OAI22_X1 U2430 ( .A1(n6364), .A2(n6691), .B1(net86719), .B2(n6359), .ZN(
        n2709) );
  OAI22_X1 U2431 ( .A1(n6364), .A2(n6694), .B1(net86720), .B2(n6359), .ZN(
        n2710) );
  OAI22_X1 U2432 ( .A1(n6364), .A2(n6697), .B1(net86721), .B2(n6359), .ZN(
        n2711) );
  OAI22_X1 U2433 ( .A1(n6364), .A2(n6700), .B1(net86722), .B2(n6359), .ZN(
        n2712) );
  OAI22_X1 U2434 ( .A1(n6378), .A2(n6629), .B1(n4294), .B2(n6377), .ZN(n2753)
         );
  OAI22_X1 U2435 ( .A1(n6378), .A2(n6634), .B1(n4096), .B2(n6377), .ZN(n2754)
         );
  OAI22_X1 U2436 ( .A1(n6378), .A2(n6637), .B1(n3898), .B2(n6377), .ZN(n2755)
         );
  OAI22_X1 U2437 ( .A1(n6378), .A2(n6640), .B1(n3844), .B2(n6377), .ZN(n2756)
         );
  OAI22_X1 U2438 ( .A1(n6378), .A2(n6643), .B1(n3826), .B2(n6377), .ZN(n2757)
         );
  OAI22_X1 U2439 ( .A1(n6379), .A2(n6646), .B1(n3808), .B2(n6377), .ZN(n2758)
         );
  OAI22_X1 U2440 ( .A1(n6379), .A2(n6649), .B1(n3790), .B2(n6377), .ZN(n2759)
         );
  OAI22_X1 U2441 ( .A1(n6379), .A2(n6652), .B1(n3772), .B2(n6377), .ZN(n2760)
         );
  OAI22_X1 U2442 ( .A1(n6379), .A2(n6655), .B1(n3754), .B2(n6377), .ZN(n2761)
         );
  OAI22_X1 U2443 ( .A1(n6379), .A2(n6658), .B1(n3736), .B2(n6377), .ZN(n2762)
         );
  OAI22_X1 U2444 ( .A1(n6380), .A2(n6661), .B1(n4276), .B2(n6377), .ZN(n2763)
         );
  OAI22_X1 U2445 ( .A1(n6380), .A2(n6664), .B1(n4258), .B2(n6377), .ZN(n2764)
         );
  OAI22_X1 U2446 ( .A1(n6380), .A2(n6667), .B1(n4240), .B2(n2338), .ZN(n2765)
         );
  OAI22_X1 U2447 ( .A1(n6380), .A2(n6670), .B1(n4222), .B2(n2338), .ZN(n2766)
         );
  OAI22_X1 U2448 ( .A1(n6380), .A2(n6673), .B1(n4204), .B2(n2338), .ZN(n2767)
         );
  OAI22_X1 U2449 ( .A1(n6381), .A2(n6676), .B1(n4186), .B2(n2338), .ZN(n2768)
         );
  OAI22_X1 U2450 ( .A1(n6381), .A2(n6679), .B1(n4168), .B2(n2338), .ZN(n2769)
         );
  OAI22_X1 U2451 ( .A1(n6381), .A2(n6682), .B1(n4150), .B2(n2338), .ZN(n2770)
         );
  OAI22_X1 U2452 ( .A1(n6381), .A2(n6685), .B1(n4132), .B2(n2338), .ZN(n2771)
         );
  OAI22_X1 U2453 ( .A1(n6381), .A2(n6688), .B1(n4114), .B2(n2338), .ZN(n2772)
         );
  OAI22_X1 U2454 ( .A1(n6382), .A2(n6691), .B1(n4078), .B2(n6377), .ZN(n2773)
         );
  OAI22_X1 U2455 ( .A1(n6382), .A2(n6694), .B1(n4060), .B2(n6377), .ZN(n2774)
         );
  OAI22_X1 U2456 ( .A1(n6382), .A2(n6697), .B1(n4042), .B2(n6377), .ZN(n2775)
         );
  OAI22_X1 U2457 ( .A1(n6382), .A2(n6700), .B1(n4024), .B2(n6377), .ZN(n2776)
         );
  OAI22_X1 U2458 ( .A1(n6387), .A2(n6629), .B1(net86731), .B2(n6386), .ZN(
        n2785) );
  OAI22_X1 U2459 ( .A1(n6387), .A2(n6634), .B1(net86732), .B2(n6386), .ZN(
        n2786) );
  OAI22_X1 U2460 ( .A1(n6387), .A2(n6637), .B1(net86733), .B2(n6386), .ZN(
        n2787) );
  OAI22_X1 U2461 ( .A1(n6387), .A2(n6640), .B1(net86734), .B2(n6386), .ZN(
        n2788) );
  OAI22_X1 U2462 ( .A1(n6387), .A2(n6643), .B1(net86735), .B2(n6386), .ZN(
        n2789) );
  OAI22_X1 U2463 ( .A1(n6388), .A2(n6646), .B1(net86736), .B2(n6386), .ZN(
        n2790) );
  OAI22_X1 U2464 ( .A1(n6388), .A2(n6649), .B1(net86737), .B2(n6386), .ZN(
        n2791) );
  OAI22_X1 U2465 ( .A1(n6388), .A2(n6652), .B1(net86738), .B2(n6386), .ZN(
        n2792) );
  OAI22_X1 U2466 ( .A1(n6388), .A2(n6655), .B1(net86739), .B2(n6386), .ZN(
        n2793) );
  OAI22_X1 U2467 ( .A1(n6388), .A2(n6658), .B1(net86740), .B2(n6386), .ZN(
        n2794) );
  OAI22_X1 U2468 ( .A1(n6389), .A2(n6661), .B1(net86741), .B2(n6386), .ZN(
        n2795) );
  OAI22_X1 U2469 ( .A1(n6389), .A2(n6664), .B1(net86742), .B2(n6386), .ZN(
        n2796) );
  OAI22_X1 U2470 ( .A1(n6389), .A2(n6667), .B1(net86743), .B2(n2336), .ZN(
        n2797) );
  OAI22_X1 U2471 ( .A1(n6389), .A2(n6670), .B1(net86744), .B2(n2336), .ZN(
        n2798) );
  OAI22_X1 U2472 ( .A1(n6389), .A2(n6673), .B1(net86745), .B2(n2336), .ZN(
        n2799) );
  OAI22_X1 U2473 ( .A1(n6390), .A2(n6676), .B1(net86746), .B2(n2336), .ZN(
        n2800) );
  OAI22_X1 U2474 ( .A1(n6390), .A2(n6679), .B1(net86747), .B2(n2336), .ZN(
        n2801) );
  OAI22_X1 U2475 ( .A1(n6390), .A2(n6682), .B1(net86748), .B2(n2336), .ZN(
        n2802) );
  OAI22_X1 U2476 ( .A1(n6390), .A2(n6685), .B1(net86749), .B2(n2336), .ZN(
        n2803) );
  OAI22_X1 U2477 ( .A1(n6390), .A2(n6688), .B1(net86750), .B2(n2336), .ZN(
        n2804) );
  OAI22_X1 U2478 ( .A1(n6391), .A2(n6691), .B1(net86751), .B2(n6386), .ZN(
        n2805) );
  OAI22_X1 U2479 ( .A1(n6391), .A2(n6694), .B1(net86752), .B2(n6386), .ZN(
        n2806) );
  OAI22_X1 U2480 ( .A1(n6391), .A2(n6697), .B1(net86753), .B2(n6386), .ZN(
        n2807) );
  OAI22_X1 U2481 ( .A1(n6391), .A2(n6700), .B1(net86754), .B2(n6386), .ZN(
        n2808) );
  OAI22_X1 U2482 ( .A1(n6396), .A2(n6629), .B1(net86763), .B2(n6395), .ZN(
        n2817) );
  OAI22_X1 U2483 ( .A1(n6396), .A2(n6634), .B1(net86764), .B2(n6395), .ZN(
        n2818) );
  OAI22_X1 U2484 ( .A1(n6396), .A2(n6637), .B1(net86765), .B2(n6395), .ZN(
        n2819) );
  OAI22_X1 U2485 ( .A1(n6396), .A2(n6640), .B1(net86766), .B2(n6395), .ZN(
        n2820) );
  OAI22_X1 U2486 ( .A1(n6396), .A2(n6643), .B1(net86767), .B2(n6395), .ZN(
        n2821) );
  OAI22_X1 U2487 ( .A1(n6397), .A2(n6646), .B1(net86768), .B2(n6395), .ZN(
        n2822) );
  OAI22_X1 U2488 ( .A1(n6397), .A2(n6649), .B1(net86769), .B2(n6395), .ZN(
        n2823) );
  OAI22_X1 U2489 ( .A1(n6397), .A2(n6652), .B1(net86770), .B2(n6395), .ZN(
        n2824) );
  OAI22_X1 U2490 ( .A1(n6397), .A2(n6655), .B1(net86771), .B2(n6395), .ZN(
        n2825) );
  OAI22_X1 U2491 ( .A1(n6397), .A2(n6658), .B1(net86772), .B2(n6395), .ZN(
        n2826) );
  OAI22_X1 U2492 ( .A1(n6398), .A2(n6661), .B1(net86773), .B2(n6395), .ZN(
        n2827) );
  OAI22_X1 U2493 ( .A1(n6398), .A2(n6664), .B1(net86774), .B2(n6395), .ZN(
        n2828) );
  OAI22_X1 U2494 ( .A1(n6398), .A2(n6667), .B1(net86775), .B2(n2334), .ZN(
        n2829) );
  OAI22_X1 U2495 ( .A1(n6398), .A2(n6670), .B1(net86776), .B2(n2334), .ZN(
        n2830) );
  OAI22_X1 U2496 ( .A1(n6398), .A2(n6673), .B1(net86777), .B2(n2334), .ZN(
        n2831) );
  OAI22_X1 U2497 ( .A1(n6399), .A2(n6676), .B1(net86778), .B2(n2334), .ZN(
        n2832) );
  OAI22_X1 U2498 ( .A1(n6399), .A2(n6679), .B1(net86779), .B2(n2334), .ZN(
        n2833) );
  OAI22_X1 U2499 ( .A1(n6399), .A2(n6682), .B1(net86780), .B2(n2334), .ZN(
        n2834) );
  OAI22_X1 U2500 ( .A1(n6399), .A2(n6685), .B1(net86781), .B2(n2334), .ZN(
        n2835) );
  OAI22_X1 U2501 ( .A1(n6399), .A2(n6688), .B1(net86782), .B2(n2334), .ZN(
        n2836) );
  OAI22_X1 U2502 ( .A1(n6400), .A2(n6691), .B1(net86783), .B2(n6395), .ZN(
        n2837) );
  OAI22_X1 U2503 ( .A1(n6400), .A2(n6694), .B1(net86784), .B2(n6395), .ZN(
        n2838) );
  OAI22_X1 U2504 ( .A1(n6400), .A2(n6697), .B1(net86785), .B2(n6395), .ZN(
        n2839) );
  OAI22_X1 U2505 ( .A1(n6400), .A2(n6700), .B1(net86786), .B2(n6395), .ZN(
        n2840) );
  OAI22_X1 U2506 ( .A1(n6423), .A2(n6629), .B1(net86795), .B2(n6422), .ZN(
        n2913) );
  OAI22_X1 U2507 ( .A1(n6423), .A2(n6633), .B1(net86796), .B2(n6422), .ZN(
        n2914) );
  OAI22_X1 U2508 ( .A1(n6423), .A2(n6636), .B1(net86797), .B2(n6422), .ZN(
        n2915) );
  OAI22_X1 U2509 ( .A1(n6423), .A2(n6639), .B1(net86798), .B2(n6422), .ZN(
        n2916) );
  OAI22_X1 U2510 ( .A1(n6423), .A2(n6642), .B1(net86799), .B2(n6422), .ZN(
        n2917) );
  OAI22_X1 U2511 ( .A1(n6424), .A2(n6645), .B1(net86800), .B2(n6422), .ZN(
        n2918) );
  OAI22_X1 U2512 ( .A1(n6424), .A2(n6648), .B1(net86801), .B2(n6422), .ZN(
        n2919) );
  OAI22_X1 U2513 ( .A1(n6424), .A2(n6651), .B1(net86802), .B2(n6422), .ZN(
        n2920) );
  OAI22_X1 U2514 ( .A1(n6424), .A2(n6654), .B1(net86803), .B2(n6422), .ZN(
        n2921) );
  OAI22_X1 U2515 ( .A1(n6424), .A2(n6657), .B1(net86804), .B2(n6422), .ZN(
        n2922) );
  OAI22_X1 U2516 ( .A1(n6425), .A2(n6660), .B1(net86805), .B2(n6422), .ZN(
        n2923) );
  OAI22_X1 U2517 ( .A1(n6425), .A2(n6663), .B1(net86806), .B2(n6422), .ZN(
        n2924) );
  OAI22_X1 U2518 ( .A1(n6425), .A2(n6666), .B1(net86807), .B2(n2277), .ZN(
        n2925) );
  OAI22_X1 U2519 ( .A1(n6425), .A2(n6669), .B1(net86808), .B2(n2277), .ZN(
        n2926) );
  OAI22_X1 U2520 ( .A1(n6425), .A2(n6672), .B1(net86809), .B2(n2277), .ZN(
        n2927) );
  OAI22_X1 U2521 ( .A1(n6426), .A2(n6675), .B1(net86810), .B2(n2277), .ZN(
        n2928) );
  OAI22_X1 U2522 ( .A1(n6426), .A2(n6678), .B1(net86811), .B2(n2277), .ZN(
        n2929) );
  OAI22_X1 U2523 ( .A1(n6426), .A2(n6681), .B1(net86812), .B2(n2277), .ZN(
        n2930) );
  OAI22_X1 U2524 ( .A1(n6426), .A2(n6684), .B1(net86813), .B2(n2277), .ZN(
        n2931) );
  OAI22_X1 U2525 ( .A1(n6426), .A2(n6687), .B1(net86814), .B2(n2277), .ZN(
        n2932) );
  OAI22_X1 U2526 ( .A1(n6427), .A2(n6690), .B1(net86815), .B2(n6422), .ZN(
        n2933) );
  OAI22_X1 U2527 ( .A1(n6427), .A2(n6693), .B1(net86816), .B2(n6422), .ZN(
        n2934) );
  OAI22_X1 U2528 ( .A1(n6427), .A2(n6696), .B1(net86817), .B2(n6422), .ZN(
        n2935) );
  OAI22_X1 U2529 ( .A1(n6427), .A2(n6699), .B1(net86818), .B2(n6422), .ZN(
        n2936) );
  OAI22_X1 U2530 ( .A1(n6432), .A2(n6629), .B1(net86827), .B2(n6431), .ZN(
        n2945) );
  OAI22_X1 U2531 ( .A1(n6432), .A2(n6633), .B1(net86828), .B2(n6431), .ZN(
        n2946) );
  OAI22_X1 U2532 ( .A1(n6432), .A2(n6636), .B1(net86829), .B2(n6431), .ZN(
        n2947) );
  OAI22_X1 U2533 ( .A1(n6432), .A2(n6639), .B1(net86830), .B2(n6431), .ZN(
        n2948) );
  OAI22_X1 U2534 ( .A1(n6432), .A2(n6642), .B1(net86831), .B2(n6431), .ZN(
        n2949) );
  OAI22_X1 U2535 ( .A1(n6433), .A2(n6645), .B1(net86832), .B2(n6431), .ZN(
        n2950) );
  OAI22_X1 U2536 ( .A1(n6433), .A2(n6648), .B1(net86833), .B2(n6431), .ZN(
        n2951) );
  OAI22_X1 U2537 ( .A1(n6433), .A2(n6651), .B1(net86834), .B2(n6431), .ZN(
        n2952) );
  OAI22_X1 U2538 ( .A1(n6433), .A2(n6654), .B1(net86835), .B2(n6431), .ZN(
        n2953) );
  OAI22_X1 U2539 ( .A1(n6433), .A2(n6657), .B1(net86836), .B2(n6431), .ZN(
        n2954) );
  OAI22_X1 U2540 ( .A1(n6434), .A2(n6660), .B1(net86837), .B2(n6431), .ZN(
        n2955) );
  OAI22_X1 U2541 ( .A1(n6434), .A2(n6663), .B1(net86838), .B2(n6431), .ZN(
        n2956) );
  OAI22_X1 U2542 ( .A1(n6434), .A2(n6666), .B1(net86839), .B2(n2275), .ZN(
        n2957) );
  OAI22_X1 U2543 ( .A1(n6434), .A2(n6669), .B1(net86840), .B2(n2275), .ZN(
        n2958) );
  OAI22_X1 U2544 ( .A1(n6434), .A2(n6672), .B1(net86841), .B2(n2275), .ZN(
        n2959) );
  OAI22_X1 U2545 ( .A1(n6435), .A2(n6675), .B1(net86842), .B2(n2275), .ZN(
        n2960) );
  OAI22_X1 U2546 ( .A1(n6435), .A2(n6678), .B1(net86843), .B2(n2275), .ZN(
        n2961) );
  OAI22_X1 U2547 ( .A1(n6435), .A2(n6681), .B1(net86844), .B2(n2275), .ZN(
        n2962) );
  OAI22_X1 U2548 ( .A1(n6435), .A2(n6684), .B1(net86845), .B2(n2275), .ZN(
        n2963) );
  OAI22_X1 U2549 ( .A1(n6435), .A2(n6687), .B1(net86846), .B2(n2275), .ZN(
        n2964) );
  OAI22_X1 U2550 ( .A1(n6436), .A2(n6690), .B1(net86847), .B2(n6431), .ZN(
        n2965) );
  OAI22_X1 U2551 ( .A1(n6436), .A2(n6693), .B1(net86848), .B2(n6431), .ZN(
        n2966) );
  OAI22_X1 U2552 ( .A1(n6436), .A2(n6696), .B1(net86849), .B2(n6431), .ZN(
        n2967) );
  OAI22_X1 U2553 ( .A1(n6436), .A2(n6699), .B1(net86850), .B2(n6431), .ZN(
        n2968) );
  OAI22_X1 U2554 ( .A1(n6459), .A2(n6630), .B1(net86859), .B2(n6458), .ZN(
        n3041) );
  OAI22_X1 U2555 ( .A1(n6459), .A2(n6633), .B1(net86860), .B2(n6458), .ZN(
        n3042) );
  OAI22_X1 U2556 ( .A1(n6459), .A2(n6636), .B1(net86861), .B2(n6458), .ZN(
        n3043) );
  OAI22_X1 U2557 ( .A1(n6459), .A2(n6639), .B1(net86862), .B2(n6458), .ZN(
        n3044) );
  OAI22_X1 U2558 ( .A1(n6459), .A2(n6642), .B1(net86863), .B2(n6458), .ZN(
        n3045) );
  OAI22_X1 U2559 ( .A1(n6460), .A2(n6645), .B1(net86864), .B2(n6458), .ZN(
        n3046) );
  OAI22_X1 U2560 ( .A1(n6460), .A2(n6648), .B1(net86865), .B2(n6458), .ZN(
        n3047) );
  OAI22_X1 U2561 ( .A1(n6460), .A2(n6651), .B1(net86866), .B2(n6458), .ZN(
        n3048) );
  OAI22_X1 U2562 ( .A1(n6460), .A2(n6654), .B1(net86867), .B2(n6458), .ZN(
        n3049) );
  OAI22_X1 U2563 ( .A1(n6460), .A2(n6657), .B1(net86868), .B2(n6458), .ZN(
        n3050) );
  OAI22_X1 U2564 ( .A1(n6461), .A2(n6660), .B1(net86869), .B2(n6458), .ZN(
        n3051) );
  OAI22_X1 U2565 ( .A1(n6461), .A2(n6663), .B1(net86870), .B2(n6458), .ZN(
        n3052) );
  OAI22_X1 U2566 ( .A1(n6461), .A2(n6666), .B1(net86871), .B2(n2217), .ZN(
        n3053) );
  OAI22_X1 U2567 ( .A1(n6461), .A2(n6669), .B1(net86872), .B2(n2217), .ZN(
        n3054) );
  OAI22_X1 U2568 ( .A1(n6461), .A2(n6672), .B1(net86873), .B2(n2217), .ZN(
        n3055) );
  OAI22_X1 U2569 ( .A1(n6462), .A2(n6675), .B1(net86874), .B2(n2217), .ZN(
        n3056) );
  OAI22_X1 U2570 ( .A1(n6462), .A2(n6678), .B1(net86875), .B2(n2217), .ZN(
        n3057) );
  OAI22_X1 U2571 ( .A1(n6462), .A2(n6681), .B1(net86876), .B2(n2217), .ZN(
        n3058) );
  OAI22_X1 U2572 ( .A1(n6462), .A2(n6684), .B1(net86877), .B2(n2217), .ZN(
        n3059) );
  OAI22_X1 U2573 ( .A1(n6462), .A2(n6687), .B1(net86878), .B2(n2217), .ZN(
        n3060) );
  OAI22_X1 U2574 ( .A1(n6463), .A2(n6690), .B1(net86879), .B2(n6458), .ZN(
        n3061) );
  OAI22_X1 U2575 ( .A1(n6463), .A2(n6693), .B1(net86880), .B2(n6458), .ZN(
        n3062) );
  OAI22_X1 U2576 ( .A1(n6463), .A2(n6696), .B1(net86881), .B2(n6458), .ZN(
        n3063) );
  OAI22_X1 U2577 ( .A1(n6463), .A2(n6699), .B1(net86882), .B2(n6458), .ZN(
        n3064) );
  OAI22_X1 U2578 ( .A1(n6468), .A2(n6630), .B1(net86891), .B2(n6467), .ZN(
        n3073) );
  OAI22_X1 U2579 ( .A1(n6468), .A2(n6633), .B1(net86892), .B2(n6467), .ZN(
        n3074) );
  OAI22_X1 U2580 ( .A1(n6468), .A2(n6636), .B1(net86893), .B2(n6467), .ZN(
        n3075) );
  OAI22_X1 U2581 ( .A1(n6468), .A2(n6639), .B1(net86894), .B2(n6467), .ZN(
        n3076) );
  OAI22_X1 U2582 ( .A1(n6468), .A2(n6642), .B1(net86895), .B2(n6467), .ZN(
        n3077) );
  OAI22_X1 U2583 ( .A1(n6469), .A2(n6645), .B1(net86896), .B2(n6467), .ZN(
        n3078) );
  OAI22_X1 U2584 ( .A1(n6469), .A2(n6648), .B1(net86897), .B2(n6467), .ZN(
        n3079) );
  OAI22_X1 U2585 ( .A1(n6469), .A2(n6651), .B1(net86898), .B2(n6467), .ZN(
        n3080) );
  OAI22_X1 U2586 ( .A1(n6469), .A2(n6654), .B1(net86899), .B2(n6467), .ZN(
        n3081) );
  OAI22_X1 U2587 ( .A1(n6469), .A2(n6657), .B1(net86900), .B2(n6467), .ZN(
        n3082) );
  OAI22_X1 U2588 ( .A1(n6470), .A2(n6660), .B1(net86901), .B2(n6467), .ZN(
        n3083) );
  OAI22_X1 U2589 ( .A1(n6470), .A2(n6663), .B1(net86902), .B2(n6467), .ZN(
        n3084) );
  OAI22_X1 U2590 ( .A1(n6470), .A2(n6666), .B1(net86903), .B2(n2215), .ZN(
        n3085) );
  OAI22_X1 U2591 ( .A1(n6470), .A2(n6669), .B1(net86904), .B2(n2215), .ZN(
        n3086) );
  OAI22_X1 U2592 ( .A1(n6470), .A2(n6672), .B1(net86905), .B2(n2215), .ZN(
        n3087) );
  OAI22_X1 U2593 ( .A1(n6471), .A2(n6675), .B1(net86906), .B2(n2215), .ZN(
        n3088) );
  OAI22_X1 U2594 ( .A1(n6471), .A2(n6678), .B1(net86907), .B2(n2215), .ZN(
        n3089) );
  OAI22_X1 U2595 ( .A1(n6471), .A2(n6681), .B1(net86908), .B2(n2215), .ZN(
        n3090) );
  OAI22_X1 U2596 ( .A1(n6471), .A2(n6684), .B1(net86909), .B2(n2215), .ZN(
        n3091) );
  OAI22_X1 U2597 ( .A1(n6471), .A2(n6687), .B1(net86910), .B2(n2215), .ZN(
        n3092) );
  OAI22_X1 U2598 ( .A1(n6472), .A2(n6690), .B1(net86911), .B2(n6467), .ZN(
        n3093) );
  OAI22_X1 U2599 ( .A1(n6472), .A2(n6693), .B1(net86912), .B2(n6467), .ZN(
        n3094) );
  OAI22_X1 U2600 ( .A1(n6472), .A2(n6696), .B1(net86913), .B2(n6467), .ZN(
        n3095) );
  OAI22_X1 U2601 ( .A1(n6472), .A2(n6699), .B1(net86914), .B2(n6467), .ZN(
        n3096) );
  OAI22_X1 U2602 ( .A1(n6495), .A2(n6630), .B1(net86923), .B2(n6494), .ZN(
        n3169) );
  OAI22_X1 U2603 ( .A1(n6495), .A2(n6633), .B1(net86924), .B2(n6494), .ZN(
        n3170) );
  OAI22_X1 U2604 ( .A1(n6495), .A2(n6636), .B1(net86925), .B2(n6494), .ZN(
        n3171) );
  OAI22_X1 U2605 ( .A1(n6495), .A2(n6639), .B1(net86926), .B2(n6494), .ZN(
        n3172) );
  OAI22_X1 U2606 ( .A1(n6495), .A2(n6642), .B1(net86927), .B2(n6494), .ZN(
        n3173) );
  OAI22_X1 U2607 ( .A1(n6496), .A2(n6645), .B1(net86928), .B2(n6494), .ZN(
        n3174) );
  OAI22_X1 U2608 ( .A1(n6496), .A2(n6648), .B1(net86929), .B2(n6494), .ZN(
        n3175) );
  OAI22_X1 U2609 ( .A1(n6496), .A2(n6651), .B1(net86930), .B2(n6494), .ZN(
        n3176) );
  OAI22_X1 U2610 ( .A1(n6496), .A2(n6654), .B1(net86931), .B2(n6494), .ZN(
        n3177) );
  OAI22_X1 U2611 ( .A1(n6496), .A2(n6657), .B1(net86932), .B2(n6494), .ZN(
        n3178) );
  OAI22_X1 U2612 ( .A1(n6497), .A2(n6660), .B1(net86933), .B2(n6494), .ZN(
        n3179) );
  OAI22_X1 U2613 ( .A1(n6497), .A2(n6663), .B1(net86934), .B2(n6494), .ZN(
        n3180) );
  OAI22_X1 U2614 ( .A1(n6497), .A2(n6666), .B1(net86935), .B2(n2157), .ZN(
        n3181) );
  OAI22_X1 U2615 ( .A1(n6497), .A2(n6669), .B1(net86936), .B2(n2157), .ZN(
        n3182) );
  OAI22_X1 U2616 ( .A1(n6497), .A2(n6672), .B1(net86937), .B2(n2157), .ZN(
        n3183) );
  OAI22_X1 U2617 ( .A1(n6498), .A2(n6675), .B1(net86938), .B2(n2157), .ZN(
        n3184) );
  OAI22_X1 U2618 ( .A1(n6498), .A2(n6678), .B1(net86939), .B2(n2157), .ZN(
        n3185) );
  OAI22_X1 U2619 ( .A1(n6498), .A2(n6681), .B1(net86940), .B2(n2157), .ZN(
        n3186) );
  OAI22_X1 U2620 ( .A1(n6498), .A2(n6684), .B1(net86941), .B2(n2157), .ZN(
        n3187) );
  OAI22_X1 U2621 ( .A1(n6498), .A2(n6687), .B1(net86942), .B2(n2157), .ZN(
        n3188) );
  OAI22_X1 U2622 ( .A1(n6499), .A2(n6690), .B1(net86943), .B2(n6494), .ZN(
        n3189) );
  OAI22_X1 U2623 ( .A1(n6499), .A2(n6693), .B1(net86944), .B2(n6494), .ZN(
        n3190) );
  OAI22_X1 U2624 ( .A1(n6499), .A2(n6696), .B1(net86945), .B2(n6494), .ZN(
        n3191) );
  OAI22_X1 U2625 ( .A1(n6499), .A2(n6699), .B1(net86946), .B2(n6494), .ZN(
        n3192) );
  OAI22_X1 U2626 ( .A1(n6504), .A2(n6630), .B1(net86955), .B2(n6503), .ZN(
        n3201) );
  OAI22_X1 U2627 ( .A1(n6504), .A2(n6633), .B1(net86956), .B2(n6503), .ZN(
        n3202) );
  OAI22_X1 U2628 ( .A1(n6504), .A2(n6636), .B1(net86957), .B2(n6503), .ZN(
        n3203) );
  OAI22_X1 U2629 ( .A1(n6504), .A2(n6639), .B1(net86958), .B2(n6503), .ZN(
        n3204) );
  OAI22_X1 U2630 ( .A1(n6504), .A2(n6642), .B1(net86959), .B2(n6503), .ZN(
        n3205) );
  OAI22_X1 U2631 ( .A1(n6505), .A2(n6645), .B1(net86960), .B2(n6503), .ZN(
        n3206) );
  OAI22_X1 U2632 ( .A1(n6505), .A2(n6648), .B1(net86961), .B2(n6503), .ZN(
        n3207) );
  OAI22_X1 U2633 ( .A1(n6505), .A2(n6651), .B1(net86962), .B2(n6503), .ZN(
        n3208) );
  OAI22_X1 U2634 ( .A1(n6505), .A2(n6654), .B1(net86963), .B2(n6503), .ZN(
        n3209) );
  OAI22_X1 U2635 ( .A1(n6505), .A2(n6657), .B1(net86964), .B2(n6503), .ZN(
        n3210) );
  OAI22_X1 U2636 ( .A1(n6506), .A2(n6660), .B1(net86965), .B2(n6503), .ZN(
        n3211) );
  OAI22_X1 U2637 ( .A1(n6506), .A2(n6663), .B1(net86966), .B2(n6503), .ZN(
        n3212) );
  OAI22_X1 U2638 ( .A1(n6506), .A2(n6666), .B1(net86967), .B2(n2155), .ZN(
        n3213) );
  OAI22_X1 U2639 ( .A1(n6506), .A2(n6669), .B1(net86968), .B2(n2155), .ZN(
        n3214) );
  OAI22_X1 U2640 ( .A1(n6506), .A2(n6672), .B1(net86969), .B2(n2155), .ZN(
        n3215) );
  OAI22_X1 U2641 ( .A1(n6507), .A2(n6675), .B1(net86970), .B2(n2155), .ZN(
        n3216) );
  OAI22_X1 U2642 ( .A1(n6507), .A2(n6678), .B1(net86971), .B2(n2155), .ZN(
        n3217) );
  OAI22_X1 U2643 ( .A1(n6507), .A2(n6681), .B1(net86972), .B2(n2155), .ZN(
        n3218) );
  OAI22_X1 U2644 ( .A1(n6507), .A2(n6684), .B1(net86973), .B2(n2155), .ZN(
        n3219) );
  OAI22_X1 U2645 ( .A1(n6507), .A2(n6687), .B1(net86974), .B2(n2155), .ZN(
        n3220) );
  OAI22_X1 U2646 ( .A1(n6508), .A2(n6690), .B1(net86975), .B2(n6503), .ZN(
        n3221) );
  OAI22_X1 U2647 ( .A1(n6508), .A2(n6693), .B1(net86976), .B2(n6503), .ZN(
        n3222) );
  OAI22_X1 U2648 ( .A1(n6508), .A2(n6696), .B1(net86977), .B2(n6503), .ZN(
        n3223) );
  OAI22_X1 U2649 ( .A1(n6508), .A2(n6699), .B1(net86978), .B2(n6503), .ZN(
        n3224) );
  OAI22_X1 U2650 ( .A1(n6531), .A2(n6630), .B1(net86987), .B2(n6530), .ZN(
        n3297) );
  OAI22_X1 U2651 ( .A1(n6531), .A2(n6632), .B1(net86988), .B2(n6530), .ZN(
        n3298) );
  OAI22_X1 U2652 ( .A1(n6531), .A2(n6635), .B1(net86989), .B2(n6530), .ZN(
        n3299) );
  OAI22_X1 U2653 ( .A1(n6531), .A2(n6638), .B1(net86990), .B2(n6530), .ZN(
        n3300) );
  OAI22_X1 U2654 ( .A1(n6531), .A2(n6641), .B1(net86991), .B2(n6530), .ZN(
        n3301) );
  OAI22_X1 U2655 ( .A1(n6532), .A2(n6644), .B1(net86992), .B2(n6530), .ZN(
        n3302) );
  OAI22_X1 U2656 ( .A1(n6532), .A2(n6647), .B1(net86993), .B2(n6530), .ZN(
        n3303) );
  OAI22_X1 U2657 ( .A1(n6532), .A2(n6650), .B1(net86994), .B2(n6530), .ZN(
        n3304) );
  OAI22_X1 U2658 ( .A1(n6532), .A2(n6653), .B1(net86995), .B2(n6530), .ZN(
        n3305) );
  OAI22_X1 U2659 ( .A1(n6532), .A2(n6656), .B1(net86996), .B2(n6530), .ZN(
        n3306) );
  OAI22_X1 U2660 ( .A1(n6533), .A2(n6659), .B1(net86997), .B2(n6530), .ZN(
        n3307) );
  OAI22_X1 U2661 ( .A1(n6533), .A2(n6662), .B1(net86998), .B2(n6530), .ZN(
        n3308) );
  OAI22_X1 U2662 ( .A1(n6533), .A2(n6665), .B1(net86999), .B2(n2098), .ZN(
        n3309) );
  OAI22_X1 U2663 ( .A1(n6533), .A2(n6668), .B1(net87000), .B2(n2098), .ZN(
        n3310) );
  OAI22_X1 U2664 ( .A1(n6533), .A2(n6671), .B1(net87001), .B2(n2098), .ZN(
        n3311) );
  OAI22_X1 U2665 ( .A1(n6534), .A2(n6674), .B1(net87002), .B2(n2098), .ZN(
        n3312) );
  OAI22_X1 U2666 ( .A1(n6534), .A2(n6677), .B1(net87003), .B2(n2098), .ZN(
        n3313) );
  OAI22_X1 U2667 ( .A1(n6534), .A2(n6680), .B1(net87004), .B2(n2098), .ZN(
        n3314) );
  OAI22_X1 U2668 ( .A1(n6534), .A2(n6683), .B1(net87005), .B2(n2098), .ZN(
        n3315) );
  OAI22_X1 U2669 ( .A1(n6534), .A2(n6686), .B1(net87006), .B2(n2098), .ZN(
        n3316) );
  OAI22_X1 U2670 ( .A1(n6535), .A2(n6689), .B1(net87007), .B2(n6530), .ZN(
        n3317) );
  OAI22_X1 U2671 ( .A1(n6535), .A2(n6692), .B1(net87008), .B2(n6530), .ZN(
        n3318) );
  OAI22_X1 U2672 ( .A1(n6535), .A2(n6695), .B1(net87009), .B2(n6530), .ZN(
        n3319) );
  OAI22_X1 U2673 ( .A1(n6535), .A2(n6698), .B1(net87010), .B2(n6530), .ZN(
        n3320) );
  OAI22_X1 U2674 ( .A1(n6540), .A2(n6630), .B1(net87019), .B2(n6539), .ZN(
        n3329) );
  OAI22_X1 U2675 ( .A1(n6540), .A2(n6632), .B1(net87020), .B2(n6539), .ZN(
        n3330) );
  OAI22_X1 U2676 ( .A1(n6540), .A2(n6635), .B1(net87021), .B2(n6539), .ZN(
        n3331) );
  OAI22_X1 U2677 ( .A1(n6540), .A2(n6638), .B1(net87022), .B2(n6539), .ZN(
        n3332) );
  OAI22_X1 U2678 ( .A1(n6540), .A2(n6641), .B1(net87023), .B2(n6539), .ZN(
        n3333) );
  OAI22_X1 U2679 ( .A1(n6541), .A2(n6644), .B1(net87024), .B2(n6539), .ZN(
        n3334) );
  OAI22_X1 U2680 ( .A1(n6541), .A2(n6647), .B1(net87025), .B2(n6539), .ZN(
        n3335) );
  OAI22_X1 U2681 ( .A1(n6541), .A2(n6650), .B1(net87026), .B2(n6539), .ZN(
        n3336) );
  OAI22_X1 U2682 ( .A1(n6541), .A2(n6653), .B1(net87027), .B2(n6539), .ZN(
        n3337) );
  OAI22_X1 U2683 ( .A1(n6541), .A2(n6656), .B1(net87028), .B2(n6539), .ZN(
        n3338) );
  OAI22_X1 U2684 ( .A1(n6542), .A2(n6659), .B1(net87029), .B2(n6539), .ZN(
        n3339) );
  OAI22_X1 U2685 ( .A1(n6542), .A2(n6662), .B1(net87030), .B2(n6539), .ZN(
        n3340) );
  OAI22_X1 U2686 ( .A1(n6542), .A2(n6665), .B1(net87031), .B2(n2096), .ZN(
        n3341) );
  OAI22_X1 U2687 ( .A1(n6542), .A2(n6668), .B1(net87032), .B2(n2096), .ZN(
        n3342) );
  OAI22_X1 U2688 ( .A1(n6542), .A2(n6671), .B1(net87033), .B2(n2096), .ZN(
        n3343) );
  OAI22_X1 U2689 ( .A1(n6543), .A2(n6674), .B1(net87034), .B2(n2096), .ZN(
        n3344) );
  OAI22_X1 U2690 ( .A1(n6543), .A2(n6677), .B1(net87035), .B2(n2096), .ZN(
        n3345) );
  OAI22_X1 U2691 ( .A1(n6543), .A2(n6680), .B1(net87036), .B2(n2096), .ZN(
        n3346) );
  OAI22_X1 U2692 ( .A1(n6543), .A2(n6683), .B1(net87037), .B2(n2096), .ZN(
        n3347) );
  OAI22_X1 U2693 ( .A1(n6543), .A2(n6686), .B1(net87038), .B2(n2096), .ZN(
        n3348) );
  OAI22_X1 U2694 ( .A1(n6544), .A2(n6689), .B1(net87039), .B2(n6539), .ZN(
        n3349) );
  OAI22_X1 U2695 ( .A1(n6544), .A2(n6692), .B1(net87040), .B2(n6539), .ZN(
        n3350) );
  OAI22_X1 U2696 ( .A1(n6544), .A2(n6695), .B1(net87041), .B2(n6539), .ZN(
        n3351) );
  OAI22_X1 U2697 ( .A1(n6544), .A2(n6698), .B1(net87042), .B2(n6539), .ZN(
        n3352) );
  OAI22_X1 U2698 ( .A1(n6567), .A2(n6631), .B1(net87051), .B2(n6566), .ZN(
        n3425) );
  OAI22_X1 U2699 ( .A1(n6567), .A2(n6632), .B1(net87052), .B2(n6566), .ZN(
        n3426) );
  OAI22_X1 U2700 ( .A1(n6567), .A2(n6635), .B1(net87053), .B2(n6566), .ZN(
        n3427) );
  OAI22_X1 U2701 ( .A1(n6567), .A2(n6638), .B1(net87054), .B2(n6566), .ZN(
        n3428) );
  OAI22_X1 U2702 ( .A1(n6567), .A2(n6641), .B1(net87055), .B2(n6566), .ZN(
        n3429) );
  OAI22_X1 U2703 ( .A1(n6568), .A2(n6644), .B1(net87056), .B2(n6566), .ZN(
        n3430) );
  OAI22_X1 U2704 ( .A1(n6568), .A2(n6647), .B1(net87057), .B2(n6566), .ZN(
        n3431) );
  OAI22_X1 U2705 ( .A1(n6568), .A2(n6650), .B1(net87058), .B2(n6566), .ZN(
        n3432) );
  OAI22_X1 U2706 ( .A1(n6568), .A2(n6653), .B1(net87059), .B2(n6566), .ZN(
        n3433) );
  OAI22_X1 U2707 ( .A1(n6568), .A2(n6656), .B1(net87060), .B2(n6566), .ZN(
        n3434) );
  OAI22_X1 U2708 ( .A1(n6569), .A2(n6659), .B1(net87061), .B2(n6566), .ZN(
        n3435) );
  OAI22_X1 U2709 ( .A1(n6569), .A2(n6662), .B1(net87062), .B2(n6566), .ZN(
        n3436) );
  OAI22_X1 U2710 ( .A1(n6569), .A2(n6665), .B1(net87063), .B2(n2037), .ZN(
        n3437) );
  OAI22_X1 U2711 ( .A1(n6569), .A2(n6668), .B1(net87064), .B2(n2037), .ZN(
        n3438) );
  OAI22_X1 U2712 ( .A1(n6569), .A2(n6671), .B1(net87065), .B2(n2037), .ZN(
        n3439) );
  OAI22_X1 U2713 ( .A1(n6570), .A2(n6674), .B1(net87066), .B2(n2037), .ZN(
        n3440) );
  OAI22_X1 U2714 ( .A1(n6570), .A2(n6677), .B1(net87067), .B2(n2037), .ZN(
        n3441) );
  OAI22_X1 U2715 ( .A1(n6570), .A2(n6680), .B1(net87068), .B2(n2037), .ZN(
        n3442) );
  OAI22_X1 U2716 ( .A1(n6570), .A2(n6683), .B1(net87069), .B2(n2037), .ZN(
        n3443) );
  OAI22_X1 U2717 ( .A1(n6570), .A2(n6686), .B1(net87070), .B2(n2037), .ZN(
        n3444) );
  OAI22_X1 U2718 ( .A1(n6571), .A2(n6689), .B1(net87071), .B2(n6566), .ZN(
        n3445) );
  OAI22_X1 U2719 ( .A1(n6571), .A2(n6692), .B1(net87072), .B2(n6566), .ZN(
        n3446) );
  OAI22_X1 U2720 ( .A1(n6571), .A2(n6695), .B1(net87073), .B2(n6566), .ZN(
        n3447) );
  OAI22_X1 U2721 ( .A1(n6571), .A2(n6698), .B1(net87074), .B2(n6566), .ZN(
        n3448) );
  OAI22_X1 U2722 ( .A1(n6576), .A2(n6631), .B1(net87083), .B2(n6575), .ZN(
        n3457) );
  OAI22_X1 U2723 ( .A1(n6576), .A2(n6632), .B1(net87084), .B2(n6575), .ZN(
        n3458) );
  OAI22_X1 U2724 ( .A1(n6576), .A2(n6635), .B1(net87085), .B2(n6575), .ZN(
        n3459) );
  OAI22_X1 U2725 ( .A1(n6576), .A2(n6638), .B1(net87086), .B2(n6575), .ZN(
        n3460) );
  OAI22_X1 U2726 ( .A1(n6576), .A2(n6641), .B1(net87087), .B2(n6575), .ZN(
        n3461) );
  OAI22_X1 U2727 ( .A1(n6577), .A2(n6644), .B1(net87088), .B2(n6575), .ZN(
        n3462) );
  OAI22_X1 U2728 ( .A1(n6577), .A2(n6647), .B1(net87089), .B2(n6575), .ZN(
        n3463) );
  OAI22_X1 U2729 ( .A1(n6577), .A2(n6650), .B1(net87090), .B2(n6575), .ZN(
        n3464) );
  OAI22_X1 U2730 ( .A1(n6577), .A2(n6653), .B1(net87091), .B2(n6575), .ZN(
        n3465) );
  OAI22_X1 U2731 ( .A1(n6577), .A2(n6656), .B1(net87092), .B2(n6575), .ZN(
        n3466) );
  OAI22_X1 U2732 ( .A1(n6578), .A2(n6659), .B1(net87093), .B2(n6575), .ZN(
        n3467) );
  OAI22_X1 U2733 ( .A1(n6578), .A2(n6662), .B1(net87094), .B2(n6575), .ZN(
        n3468) );
  OAI22_X1 U2734 ( .A1(n6578), .A2(n6665), .B1(net87095), .B2(n2035), .ZN(
        n3469) );
  OAI22_X1 U2735 ( .A1(n6578), .A2(n6668), .B1(net87096), .B2(n2035), .ZN(
        n3470) );
  OAI22_X1 U2736 ( .A1(n6578), .A2(n6671), .B1(net87097), .B2(n2035), .ZN(
        n3471) );
  OAI22_X1 U2737 ( .A1(n6579), .A2(n6674), .B1(net87098), .B2(n2035), .ZN(
        n3472) );
  OAI22_X1 U2738 ( .A1(n6579), .A2(n6677), .B1(net87099), .B2(n2035), .ZN(
        n3473) );
  OAI22_X1 U2739 ( .A1(n6579), .A2(n6680), .B1(net87100), .B2(n2035), .ZN(
        n3474) );
  OAI22_X1 U2740 ( .A1(n6579), .A2(n6683), .B1(net87101), .B2(n2035), .ZN(
        n3475) );
  OAI22_X1 U2741 ( .A1(n6579), .A2(n6686), .B1(net87102), .B2(n2035), .ZN(
        n3476) );
  OAI22_X1 U2742 ( .A1(n6580), .A2(n6689), .B1(net87103), .B2(n6575), .ZN(
        n3477) );
  OAI22_X1 U2743 ( .A1(n6580), .A2(n6692), .B1(net87104), .B2(n6575), .ZN(
        n3478) );
  OAI22_X1 U2744 ( .A1(n6580), .A2(n6695), .B1(net87105), .B2(n6575), .ZN(
        n3479) );
  OAI22_X1 U2745 ( .A1(n6580), .A2(n6698), .B1(net87106), .B2(n6575), .ZN(
        n3480) );
  OAI22_X1 U2746 ( .A1(n6603), .A2(n6631), .B1(net87115), .B2(n6602), .ZN(
        n3553) );
  OAI22_X1 U2747 ( .A1(n6603), .A2(n6632), .B1(net87116), .B2(n6602), .ZN(
        n3554) );
  OAI22_X1 U2748 ( .A1(n6603), .A2(n6635), .B1(net87117), .B2(n6602), .ZN(
        n3555) );
  OAI22_X1 U2749 ( .A1(n6603), .A2(n6638), .B1(net87118), .B2(n6602), .ZN(
        n3556) );
  OAI22_X1 U2750 ( .A1(n6603), .A2(n6641), .B1(net87119), .B2(n6602), .ZN(
        n3557) );
  OAI22_X1 U2751 ( .A1(n6604), .A2(n6644), .B1(net87120), .B2(n6602), .ZN(
        n3558) );
  OAI22_X1 U2752 ( .A1(n6604), .A2(n6647), .B1(net87121), .B2(n6602), .ZN(
        n3559) );
  OAI22_X1 U2753 ( .A1(n6604), .A2(n6650), .B1(net87122), .B2(n6602), .ZN(
        n3560) );
  OAI22_X1 U2754 ( .A1(n6604), .A2(n6653), .B1(net87123), .B2(n6602), .ZN(
        n3561) );
  OAI22_X1 U2755 ( .A1(n6604), .A2(n6656), .B1(net87124), .B2(n6602), .ZN(
        n3562) );
  OAI22_X1 U2756 ( .A1(n6605), .A2(n6659), .B1(net87125), .B2(n6602), .ZN(
        n3563) );
  OAI22_X1 U2757 ( .A1(n6605), .A2(n6662), .B1(net87126), .B2(n6602), .ZN(
        n3564) );
  OAI22_X1 U2758 ( .A1(n6605), .A2(n6665), .B1(net87127), .B2(n1972), .ZN(
        n3565) );
  OAI22_X1 U2759 ( .A1(n6605), .A2(n6668), .B1(net87128), .B2(n1972), .ZN(
        n3566) );
  OAI22_X1 U2760 ( .A1(n6605), .A2(n6671), .B1(net87129), .B2(n1972), .ZN(
        n3567) );
  OAI22_X1 U2761 ( .A1(n6606), .A2(n6674), .B1(net87130), .B2(n1972), .ZN(
        n3568) );
  OAI22_X1 U2762 ( .A1(n6606), .A2(n6677), .B1(net87131), .B2(n1972), .ZN(
        n3569) );
  OAI22_X1 U2763 ( .A1(n6606), .A2(n6680), .B1(net87132), .B2(n1972), .ZN(
        n3570) );
  OAI22_X1 U2764 ( .A1(n6606), .A2(n6683), .B1(net87133), .B2(n1972), .ZN(
        n3571) );
  OAI22_X1 U2765 ( .A1(n6606), .A2(n6686), .B1(net87134), .B2(n1972), .ZN(
        n3572) );
  OAI22_X1 U2766 ( .A1(n6607), .A2(n6689), .B1(net87135), .B2(n6602), .ZN(
        n3573) );
  OAI22_X1 U2767 ( .A1(n6607), .A2(n6692), .B1(net87136), .B2(n6602), .ZN(
        n3574) );
  OAI22_X1 U2768 ( .A1(n6607), .A2(n6695), .B1(net87137), .B2(n6602), .ZN(
        n3575) );
  OAI22_X1 U2769 ( .A1(n6607), .A2(n6698), .B1(net87138), .B2(n6602), .ZN(
        n3576) );
  OAI22_X1 U2770 ( .A1(n6612), .A2(n6631), .B1(net87147), .B2(n6611), .ZN(
        n3585) );
  OAI22_X1 U2771 ( .A1(n6612), .A2(n6632), .B1(net87148), .B2(n6611), .ZN(
        n3586) );
  OAI22_X1 U2772 ( .A1(n6612), .A2(n6635), .B1(net87149), .B2(n6611), .ZN(
        n3587) );
  OAI22_X1 U2773 ( .A1(n6612), .A2(n6638), .B1(net87150), .B2(n6611), .ZN(
        n3588) );
  OAI22_X1 U2774 ( .A1(n6612), .A2(n6641), .B1(net87151), .B2(n6611), .ZN(
        n3589) );
  OAI22_X1 U2775 ( .A1(n6613), .A2(n6644), .B1(net87152), .B2(n6611), .ZN(
        n3590) );
  OAI22_X1 U2776 ( .A1(n6613), .A2(n6647), .B1(net87153), .B2(n6611), .ZN(
        n3591) );
  OAI22_X1 U2777 ( .A1(n6613), .A2(n6650), .B1(net87154), .B2(n6611), .ZN(
        n3592) );
  OAI22_X1 U2778 ( .A1(n6613), .A2(n6653), .B1(net87155), .B2(n6611), .ZN(
        n3593) );
  OAI22_X1 U2779 ( .A1(n6613), .A2(n6656), .B1(net87156), .B2(n6611), .ZN(
        n3594) );
  OAI22_X1 U2780 ( .A1(n6614), .A2(n6659), .B1(net87157), .B2(n6611), .ZN(
        n3595) );
  OAI22_X1 U2781 ( .A1(n6614), .A2(n6662), .B1(net87158), .B2(n6611), .ZN(
        n3596) );
  OAI22_X1 U2782 ( .A1(n6614), .A2(n6665), .B1(net87159), .B2(n1969), .ZN(
        n3597) );
  OAI22_X1 U2783 ( .A1(n6614), .A2(n6668), .B1(net87160), .B2(n1969), .ZN(
        n3598) );
  OAI22_X1 U2784 ( .A1(n6614), .A2(n6671), .B1(net87161), .B2(n1969), .ZN(
        n3599) );
  OAI22_X1 U2785 ( .A1(n6615), .A2(n6674), .B1(net87162), .B2(n1969), .ZN(
        n3600) );
  OAI22_X1 U2786 ( .A1(n6615), .A2(n6677), .B1(net87163), .B2(n1969), .ZN(
        n3601) );
  OAI22_X1 U2787 ( .A1(n6615), .A2(n6680), .B1(net87164), .B2(n1969), .ZN(
        n3602) );
  OAI22_X1 U2788 ( .A1(n6615), .A2(n6683), .B1(net87165), .B2(n1969), .ZN(
        n3603) );
  OAI22_X1 U2789 ( .A1(n6615), .A2(n6686), .B1(net87166), .B2(n1969), .ZN(
        n3604) );
  OAI22_X1 U2790 ( .A1(n6616), .A2(n6689), .B1(net87167), .B2(n6611), .ZN(
        n3605) );
  OAI22_X1 U2791 ( .A1(n6616), .A2(n6692), .B1(net87168), .B2(n6611), .ZN(
        n3606) );
  OAI22_X1 U2792 ( .A1(n6616), .A2(n6695), .B1(net87169), .B2(n6611), .ZN(
        n3607) );
  OAI22_X1 U2793 ( .A1(n6616), .A2(n6698), .B1(net87170), .B2(n6611), .ZN(
        n3608) );
  OAI22_X1 U2794 ( .A1(n6405), .A2(n6637), .B1(n68), .B2(n2310), .ZN(n2851) );
  OAI22_X1 U2795 ( .A1(n6405), .A2(n6640), .B1(n47), .B2(n2310), .ZN(n2852) );
  OAI22_X1 U2796 ( .A1(n6405), .A2(n6643), .B1(n40), .B2(n6404), .ZN(n2853) );
  OAI22_X1 U2797 ( .A1(n6406), .A2(n6658), .B1(n5), .B2(n2310), .ZN(n2858) );
  OAI22_X1 U2798 ( .A1(n6410), .A2(n6709), .B1(n96), .B2(n6404), .ZN(n2875) );
  OAI22_X1 U2799 ( .A1(n6410), .A2(n6712), .B1(n89), .B2(n2310), .ZN(n2876) );
  OAI22_X1 U2800 ( .A1(n6410), .A2(n6715), .B1(n82), .B2(n2310), .ZN(n2877) );
  OAI22_X1 U2801 ( .A1(n6410), .A2(n6718), .B1(n75), .B2(n2310), .ZN(n2878) );
  OAI22_X1 U2802 ( .A1(n6411), .A2(n6721), .B1(n61), .B2(n6404), .ZN(n2879) );
  OAI22_X1 U2803 ( .A1(n6411), .A2(n6733), .B1(n54), .B2(n6404), .ZN(n2880) );
  OAI22_X1 U2804 ( .A1(n6450), .A2(n6636), .B1(n70), .B2(n2220), .ZN(n3011) );
  OAI22_X1 U2805 ( .A1(n6450), .A2(n6639), .B1(n49), .B2(n2220), .ZN(n3012) );
  OAI22_X1 U2806 ( .A1(n6450), .A2(n6642), .B1(n42), .B2(n6449), .ZN(n3013) );
  OAI22_X1 U2807 ( .A1(n6451), .A2(n6657), .B1(n7), .B2(n2220), .ZN(n3018) );
  OAI22_X1 U2808 ( .A1(n6455), .A2(n6708), .B1(n98), .B2(n6449), .ZN(n3035) );
  OAI22_X1 U2809 ( .A1(n6455), .A2(n6711), .B1(n91), .B2(n2220), .ZN(n3036) );
  OAI22_X1 U2810 ( .A1(n6455), .A2(n6714), .B1(n84), .B2(n2220), .ZN(n3037) );
  OAI22_X1 U2811 ( .A1(n6455), .A2(n6717), .B1(n77), .B2(n2220), .ZN(n3038) );
  OAI22_X1 U2812 ( .A1(n6456), .A2(n6720), .B1(n63), .B2(n6449), .ZN(n3039) );
  OAI22_X1 U2813 ( .A1(n6456), .A2(n6732), .B1(n56), .B2(n6449), .ZN(n3040) );
  OAI22_X1 U2814 ( .A1(n6486), .A2(n6636), .B1(n69), .B2(n2160), .ZN(n3139) );
  OAI22_X1 U2815 ( .A1(n6486), .A2(n6639), .B1(n48), .B2(n2160), .ZN(n3140) );
  OAI22_X1 U2816 ( .A1(n6486), .A2(n6642), .B1(n41), .B2(n6485), .ZN(n3141) );
  OAI22_X1 U2817 ( .A1(n6487), .A2(n6657), .B1(n6), .B2(n2160), .ZN(n3146) );
  OAI22_X1 U2818 ( .A1(n6491), .A2(n6708), .B1(n97), .B2(n6485), .ZN(n3163) );
  OAI22_X1 U2819 ( .A1(n6491), .A2(n6711), .B1(n90), .B2(n2160), .ZN(n3164) );
  OAI22_X1 U2820 ( .A1(n6491), .A2(n6714), .B1(n83), .B2(n2160), .ZN(n3165) );
  OAI22_X1 U2821 ( .A1(n6491), .A2(n6717), .B1(n76), .B2(n2160), .ZN(n3166) );
  OAI22_X1 U2822 ( .A1(n6492), .A2(n6720), .B1(n62), .B2(n6485), .ZN(n3167) );
  OAI22_X1 U2823 ( .A1(n6492), .A2(n6732), .B1(n55), .B2(n6485), .ZN(n3168) );
  OAI22_X1 U2824 ( .A1(n6513), .A2(n6636), .B1(n67), .B2(n2131), .ZN(n3235) );
  OAI22_X1 U2825 ( .A1(n6513), .A2(n6639), .B1(n46), .B2(n2131), .ZN(n3236) );
  OAI22_X1 U2826 ( .A1(n6513), .A2(n6642), .B1(n39), .B2(n6512), .ZN(n3237) );
  OAI22_X1 U2827 ( .A1(n6514), .A2(n6657), .B1(n4), .B2(n2131), .ZN(n3242) );
  OAI22_X1 U2828 ( .A1(n6518), .A2(n6708), .B1(n95), .B2(n6512), .ZN(n3259) );
  OAI22_X1 U2829 ( .A1(n6518), .A2(n6711), .B1(n88), .B2(n2131), .ZN(n3260) );
  OAI22_X1 U2830 ( .A1(n6518), .A2(n6714), .B1(n81), .B2(n2131), .ZN(n3261) );
  OAI22_X1 U2831 ( .A1(n6518), .A2(n6717), .B1(n74), .B2(n2131), .ZN(n3262) );
  OAI22_X1 U2832 ( .A1(n6519), .A2(n6720), .B1(n60), .B2(n6512), .ZN(n3263) );
  OAI22_X1 U2833 ( .A1(n6519), .A2(n6732), .B1(n53), .B2(n6512), .ZN(n3264) );
  OAI22_X1 U2834 ( .A1(n6621), .A2(n6635), .B1(n64), .B2(n1944), .ZN(n3619) );
  OAI22_X1 U2835 ( .A1(n6621), .A2(n6638), .B1(n43), .B2(n1944), .ZN(n3620) );
  OAI22_X1 U2836 ( .A1(n6622), .A2(n6653), .B1(n8), .B2(n6620), .ZN(n3625) );
  OAI22_X1 U2837 ( .A1(n6626), .A2(n6704), .B1(n99), .B2(n1944), .ZN(n3642) );
  OAI22_X1 U2838 ( .A1(n6626), .A2(n6707), .B1(n92), .B2(n6620), .ZN(n3643) );
  OAI22_X1 U2839 ( .A1(n6626), .A2(n6710), .B1(n85), .B2(n1944), .ZN(n3644) );
  OAI22_X1 U2840 ( .A1(n6626), .A2(n6713), .B1(n78), .B2(n1944), .ZN(n3645) );
  OAI22_X1 U2841 ( .A1(n6626), .A2(n6716), .B1(n71), .B2(n1944), .ZN(n3646) );
  OAI22_X1 U2842 ( .A1(n6627), .A2(n6719), .B1(n57), .B2(n1944), .ZN(n3647) );
  OAI22_X1 U2843 ( .A1(n6627), .A2(n6731), .B1(n50), .B2(n1944), .ZN(n3648) );
  OAI22_X1 U2844 ( .A1(n6585), .A2(n6635), .B1(n65), .B2(n2010), .ZN(n3491) );
  OAI22_X1 U2845 ( .A1(n6585), .A2(n6638), .B1(n44), .B2(n6584), .ZN(n3492) );
  OAI22_X1 U2846 ( .A1(n6586), .A2(n6653), .B1(n9), .B2(n6584), .ZN(n3497) );
  OAI22_X1 U2847 ( .A1(n6590), .A2(n6707), .B1(n93), .B2(n2010), .ZN(n3515) );
  OAI22_X1 U2848 ( .A1(n6590), .A2(n6710), .B1(n86), .B2(n2010), .ZN(n3516) );
  OAI22_X1 U2849 ( .A1(n6590), .A2(n6713), .B1(n79), .B2(n2010), .ZN(n3517) );
  OAI22_X1 U2850 ( .A1(n6590), .A2(n6716), .B1(n72), .B2(n2010), .ZN(n3518) );
  OAI22_X1 U2851 ( .A1(n6591), .A2(n6719), .B1(n58), .B2(n6584), .ZN(n3519) );
  OAI22_X1 U2852 ( .A1(n6591), .A2(n6731), .B1(n51), .B2(n6584), .ZN(n3520) );
  OAI22_X1 U2853 ( .A1(n6549), .A2(n6635), .B1(n66), .B2(n6548), .ZN(n3363) );
  OAI22_X1 U2854 ( .A1(n6549), .A2(n6638), .B1(n45), .B2(n6548), .ZN(n3364) );
  OAI22_X1 U2855 ( .A1(n6554), .A2(n6707), .B1(n94), .B2(n2070), .ZN(n3387) );
  OAI22_X1 U2856 ( .A1(n6554), .A2(n6710), .B1(n87), .B2(n6548), .ZN(n3388) );
  OAI22_X1 U2857 ( .A1(n6554), .A2(n6713), .B1(n80), .B2(n2070), .ZN(n3389) );
  OAI22_X1 U2858 ( .A1(n6554), .A2(n6716), .B1(n73), .B2(n6548), .ZN(n3390) );
  OAI22_X1 U2859 ( .A1(n6555), .A2(n6719), .B1(n59), .B2(n2070), .ZN(n3391) );
  OAI22_X1 U2860 ( .A1(n6555), .A2(n6731), .B1(n52), .B2(n2070), .ZN(n3392) );
  INV_X1 U2861 ( .A(RD2), .ZN(n5082) );
  INV_X1 U2862 ( .A(ADD_RD2[0]), .ZN(n5053) );
  INV_X1 U2863 ( .A(ADD_RD2[3]), .ZN(n5054) );
  NOR3_X1 U2864 ( .A1(n5720), .A2(n5710), .A3(n5721), .ZN(n5719) );
  XNOR2_X1 U2865 ( .A(n2340), .B(ADD_RD1[1]), .ZN(n5720) );
  XNOR2_X1 U2866 ( .A(ADD_WR[4]), .B(n5705), .ZN(n5721) );
  XNOR2_X1 U2867 ( .A(ADD_RD2[2]), .B(ADD_WR[2]), .ZN(n5722) );
  INV_X1 U2868 ( .A(ADD_WR[1]), .ZN(n2340) );
  INV_X1 U2869 ( .A(ADD_RD2[1]), .ZN(n5081) );
  INV_X1 U2870 ( .A(ADD_RD2[2]), .ZN(n5086) );
  AND2_X1 U2871 ( .A1(ADD_WR[4]), .A2(WR), .ZN(n2218) );
  INV_X1 U2872 ( .A(ADD_WR[2]), .ZN(n1974) );
  INV_X1 U2873 ( .A(WR), .ZN(n2158) );
  INV_X1 U2874 ( .A(ADD_WR[3]), .ZN(n1975) );
  XNOR2_X1 U2875 ( .A(ADD_RD1[3]), .B(ADD_WR[3]), .ZN(n5718) );
  XNOR2_X1 U2876 ( .A(ADD_RD2[3]), .B(ADD_WR[3]), .ZN(n5724) );
  XNOR2_X1 U2877 ( .A(ADD_WR[0]), .B(ADD_RD2[0]), .ZN(n5723) );
  XNOR2_X1 U2878 ( .A(ADD_WR[0]), .B(ADD_RD1[0]), .ZN(n5717) );
  NAND2_X1 U2879 ( .A1(ADD_WR[0]), .A2(n2340), .ZN(n1967) );
  NAND2_X1 U2880 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .ZN(n1973) );
  INV_X1 U2881 ( .A(ADD_WR[0]), .ZN(n2341) );
  INV_X1 U2882 ( .A(n5884), .ZN(n5885) );
  INV_X1 U2883 ( .A(n5884), .ZN(n5886) );
  INV_X1 U2884 ( .A(n5884), .ZN(n5887) );
  INV_X1 U2885 ( .A(n5884), .ZN(n5888) );
  INV_X1 U2886 ( .A(n5884), .ZN(n5889) );
  INV_X1 U2887 ( .A(n5884), .ZN(n5890) );
  INV_X1 U2888 ( .A(n5884), .ZN(n5891) );
  INV_X1 U2889 ( .A(n5892), .ZN(n5894) );
  INV_X1 U2890 ( .A(n5892), .ZN(n5895) );
  INV_X1 U2891 ( .A(n5893), .ZN(n5896) );
  INV_X1 U2892 ( .A(n5893), .ZN(n5897) );
  INV_X1 U2893 ( .A(n5892), .ZN(n5898) );
  INV_X1 U2894 ( .A(n5893), .ZN(n5899) );
  INV_X1 U2895 ( .A(n5135), .ZN(n5900) );
  INV_X1 U2896 ( .A(n5135), .ZN(n5901) );
  INV_X1 U2897 ( .A(n5901), .ZN(n5902) );
  INV_X1 U2898 ( .A(n5900), .ZN(n5903) );
  INV_X1 U2899 ( .A(n5901), .ZN(n5904) );
  INV_X1 U2900 ( .A(n5900), .ZN(n5905) );
  INV_X1 U2901 ( .A(n5901), .ZN(n5906) );
  INV_X1 U2902 ( .A(n5900), .ZN(n5907) );
  INV_X1 U2903 ( .A(n5136), .ZN(n5908) );
  INV_X1 U2904 ( .A(n5136), .ZN(n5909) );
  INV_X1 U2905 ( .A(n5908), .ZN(n5910) );
  INV_X1 U2906 ( .A(n5909), .ZN(n5911) );
  INV_X1 U2907 ( .A(n5908), .ZN(n5912) );
  INV_X1 U2908 ( .A(n5908), .ZN(n5913) );
  INV_X1 U2909 ( .A(n5908), .ZN(n5914) );
  INV_X1 U2910 ( .A(n5909), .ZN(n5915) );
  INV_X1 U2911 ( .A(n5916), .ZN(n5918) );
  INV_X1 U2912 ( .A(n5916), .ZN(n5919) );
  INV_X1 U2913 ( .A(n5917), .ZN(n5920) );
  INV_X1 U2914 ( .A(n5917), .ZN(n5921) );
  INV_X1 U2915 ( .A(n5917), .ZN(n5922) );
  INV_X1 U2916 ( .A(n5916), .ZN(n5923) );
  INV_X1 U2917 ( .A(n5924), .ZN(n5925) );
  INV_X1 U2918 ( .A(n5924), .ZN(n5926) );
  INV_X1 U2919 ( .A(n5924), .ZN(n5927) );
  INV_X1 U2920 ( .A(n5924), .ZN(n5928) );
  INV_X1 U2921 ( .A(n5924), .ZN(n5929) );
  INV_X1 U2922 ( .A(n5924), .ZN(n5930) );
  INV_X1 U2923 ( .A(n5924), .ZN(n5931) );
  INV_X1 U2924 ( .A(n5130), .ZN(n5932) );
  INV_X1 U2925 ( .A(n5932), .ZN(n5933) );
  INV_X1 U2926 ( .A(n5932), .ZN(n5934) );
  INV_X1 U2927 ( .A(n5932), .ZN(n5935) );
  INV_X1 U2928 ( .A(n5932), .ZN(n5936) );
  INV_X1 U2929 ( .A(n5932), .ZN(n5937) );
  INV_X1 U2930 ( .A(n5932), .ZN(n5938) );
  INV_X1 U2931 ( .A(n5932), .ZN(n5939) );
  INV_X1 U2932 ( .A(n5131), .ZN(n5940) );
  INV_X1 U2933 ( .A(n5940), .ZN(n5941) );
  INV_X1 U2934 ( .A(n5940), .ZN(n5942) );
  INV_X1 U2935 ( .A(n5940), .ZN(n5943) );
  INV_X1 U2936 ( .A(n5940), .ZN(n5944) );
  INV_X1 U2937 ( .A(n5940), .ZN(n5945) );
  INV_X1 U2938 ( .A(n5940), .ZN(n5946) );
  INV_X1 U2939 ( .A(n5940), .ZN(n5947) );
  INV_X1 U2940 ( .A(n5948), .ZN(n5950) );
  INV_X1 U2941 ( .A(n5949), .ZN(n5951) );
  INV_X1 U2942 ( .A(n5948), .ZN(n5952) );
  INV_X1 U2943 ( .A(n5948), .ZN(n5953) );
  INV_X1 U2944 ( .A(n5949), .ZN(n5954) );
  INV_X1 U2945 ( .A(n5949), .ZN(n5955) );
  INV_X1 U2946 ( .A(n5956), .ZN(n5958) );
  INV_X1 U2947 ( .A(n5957), .ZN(n5959) );
  INV_X1 U2948 ( .A(n5956), .ZN(n5960) );
  INV_X1 U2949 ( .A(n5956), .ZN(n5961) );
  INV_X1 U2950 ( .A(n5957), .ZN(n5962) );
  INV_X1 U2951 ( .A(n5957), .ZN(n5963) );
  INV_X1 U2952 ( .A(n5125), .ZN(n5964) );
  INV_X1 U2953 ( .A(n5964), .ZN(n5965) );
  INV_X1 U2954 ( .A(n5964), .ZN(n5966) );
  INV_X1 U2955 ( .A(n5964), .ZN(n5967) );
  INV_X1 U2956 ( .A(n5964), .ZN(n5968) );
  INV_X1 U2957 ( .A(n5964), .ZN(n5969) );
  INV_X1 U2958 ( .A(n5964), .ZN(n5970) );
  INV_X1 U2959 ( .A(n5964), .ZN(n5971) );
  INV_X1 U2960 ( .A(n5126), .ZN(n5972) );
  INV_X1 U2961 ( .A(n5972), .ZN(n5973) );
  INV_X1 U2962 ( .A(n5972), .ZN(n5974) );
  INV_X1 U2963 ( .A(n5972), .ZN(n5975) );
  INV_X1 U2964 ( .A(n5972), .ZN(n5976) );
  INV_X1 U2965 ( .A(n5972), .ZN(n5977) );
  INV_X1 U2966 ( .A(n5972), .ZN(n5978) );
  INV_X1 U2967 ( .A(n5972), .ZN(n5979) );
  INV_X1 U2968 ( .A(n5980), .ZN(n5982) );
  INV_X1 U2969 ( .A(n5981), .ZN(n5983) );
  INV_X1 U2970 ( .A(n5980), .ZN(n5984) );
  INV_X1 U2971 ( .A(n5980), .ZN(n5985) );
  INV_X1 U2972 ( .A(n5981), .ZN(n5986) );
  INV_X1 U2973 ( .A(n5981), .ZN(n5987) );
  INV_X1 U2974 ( .A(n5988), .ZN(n5990) );
  INV_X1 U2975 ( .A(n5989), .ZN(n5991) );
  INV_X1 U2976 ( .A(n5988), .ZN(n5992) );
  INV_X1 U2977 ( .A(n5988), .ZN(n5993) );
  INV_X1 U2978 ( .A(n5989), .ZN(n5994) );
  INV_X1 U2979 ( .A(n5989), .ZN(n5995) );
  INV_X1 U2980 ( .A(n5120), .ZN(n5996) );
  INV_X1 U2981 ( .A(n5996), .ZN(n5997) );
  INV_X1 U2982 ( .A(n5996), .ZN(n5998) );
  INV_X1 U2983 ( .A(n5996), .ZN(n5999) );
  INV_X1 U2984 ( .A(n5996), .ZN(n6000) );
  INV_X1 U2985 ( .A(n5996), .ZN(n6001) );
  INV_X1 U2986 ( .A(n5996), .ZN(n6002) );
  INV_X1 U2987 ( .A(n5996), .ZN(n6003) );
  INV_X1 U2988 ( .A(n5121), .ZN(n6004) );
  INV_X1 U2989 ( .A(n6004), .ZN(n6005) );
  INV_X1 U2990 ( .A(n6004), .ZN(n6006) );
  INV_X1 U2991 ( .A(n6004), .ZN(n6007) );
  INV_X1 U2992 ( .A(n6004), .ZN(n6008) );
  INV_X1 U2993 ( .A(n6004), .ZN(n6009) );
  INV_X1 U2994 ( .A(n6004), .ZN(n6010) );
  INV_X1 U2995 ( .A(n6004), .ZN(n6011) );
  INV_X1 U2996 ( .A(n6012), .ZN(n6014) );
  INV_X1 U2997 ( .A(n6012), .ZN(n6015) );
  INV_X1 U2998 ( .A(n6012), .ZN(n6016) );
  INV_X1 U2999 ( .A(n6013), .ZN(n6017) );
  INV_X1 U3000 ( .A(n6013), .ZN(n6018) );
  INV_X1 U3001 ( .A(n6013), .ZN(n6019) );
  INV_X1 U3002 ( .A(n6020), .ZN(n6021) );
  INV_X1 U3003 ( .A(n6020), .ZN(n6022) );
  INV_X1 U3004 ( .A(n6020), .ZN(n6023) );
  INV_X1 U3005 ( .A(n6020), .ZN(n6024) );
  INV_X1 U3006 ( .A(n6020), .ZN(n6025) );
  INV_X1 U3007 ( .A(n6020), .ZN(n6026) );
  INV_X1 U3008 ( .A(n6020), .ZN(n6027) );
  INV_X1 U3009 ( .A(n5111), .ZN(n6028) );
  INV_X1 U3010 ( .A(n5111), .ZN(n6029) );
  INV_X1 U3011 ( .A(n6029), .ZN(n6030) );
  INV_X1 U3012 ( .A(n6028), .ZN(n6031) );
  INV_X1 U3013 ( .A(n6028), .ZN(n6032) );
  INV_X1 U3014 ( .A(n6029), .ZN(n6033) );
  INV_X1 U3015 ( .A(n6029), .ZN(n6034) );
  INV_X1 U3016 ( .A(n6028), .ZN(n6035) );
  INV_X1 U3017 ( .A(n5112), .ZN(n6036) );
  INV_X1 U3018 ( .A(n6036), .ZN(n6037) );
  INV_X1 U3019 ( .A(n6036), .ZN(n6038) );
  INV_X1 U3020 ( .A(n6036), .ZN(n6039) );
  INV_X1 U3021 ( .A(n6036), .ZN(n6040) );
  INV_X1 U3022 ( .A(n6036), .ZN(n6041) );
  INV_X1 U3023 ( .A(n6036), .ZN(n6042) );
  INV_X1 U3024 ( .A(n6036), .ZN(n6043) );
  INV_X1 U3025 ( .A(n6044), .ZN(n6045) );
  INV_X1 U3026 ( .A(n6044), .ZN(n6046) );
  INV_X1 U3027 ( .A(n6044), .ZN(n6047) );
  INV_X1 U3028 ( .A(n6044), .ZN(n6048) );
  INV_X1 U3029 ( .A(n6044), .ZN(n6049) );
  INV_X1 U3030 ( .A(n6044), .ZN(n6050) );
  INV_X1 U3031 ( .A(n6044), .ZN(n6051) );
  INV_X1 U3032 ( .A(n6052), .ZN(n6053) );
  INV_X1 U3033 ( .A(n6052), .ZN(n6054) );
  INV_X1 U3034 ( .A(n6052), .ZN(n6055) );
  INV_X1 U3035 ( .A(n6052), .ZN(n6056) );
  INV_X1 U3036 ( .A(n6052), .ZN(n6057) );
  INV_X1 U3037 ( .A(n6052), .ZN(n6058) );
  INV_X1 U3038 ( .A(n6052), .ZN(n6059) );
  INV_X1 U3039 ( .A(n5106), .ZN(n6060) );
  INV_X1 U3040 ( .A(n6060), .ZN(n6061) );
  INV_X1 U3041 ( .A(n6060), .ZN(n6062) );
  INV_X1 U3042 ( .A(n6060), .ZN(n6063) );
  INV_X1 U3043 ( .A(n6060), .ZN(n6064) );
  INV_X1 U3044 ( .A(n6060), .ZN(n6065) );
  INV_X1 U3045 ( .A(n6060), .ZN(n6066) );
  INV_X1 U3046 ( .A(n6060), .ZN(n6067) );
  INV_X1 U3047 ( .A(n5107), .ZN(n6068) );
  INV_X1 U3048 ( .A(n5107), .ZN(n6069) );
  INV_X1 U3049 ( .A(n6069), .ZN(n6070) );
  INV_X1 U3050 ( .A(n6068), .ZN(n6071) );
  INV_X1 U3051 ( .A(n6068), .ZN(n6072) );
  INV_X1 U3052 ( .A(n6069), .ZN(n6073) );
  INV_X1 U3053 ( .A(n6069), .ZN(n6074) );
  INV_X1 U3054 ( .A(n6068), .ZN(n6075) );
  INV_X1 U3055 ( .A(n6076), .ZN(n6078) );
  INV_X1 U3056 ( .A(n6077), .ZN(n6079) );
  INV_X1 U3057 ( .A(n6077), .ZN(n6080) );
  INV_X1 U3058 ( .A(n6077), .ZN(n6081) );
  INV_X1 U3059 ( .A(n6076), .ZN(n6082) );
  INV_X1 U3060 ( .A(n6077), .ZN(n6083) );
  INV_X1 U3061 ( .A(n6084), .ZN(n6086) );
  INV_X1 U3062 ( .A(n6084), .ZN(n6087) );
  INV_X1 U3063 ( .A(n6085), .ZN(n6088) );
  INV_X1 U3064 ( .A(n6084), .ZN(n6089) );
  INV_X1 U3065 ( .A(n6085), .ZN(n6090) );
  INV_X1 U3066 ( .A(n6085), .ZN(n6091) );
  INV_X1 U3067 ( .A(n6096), .ZN(n6097) );
  INV_X1 U3068 ( .A(n6096), .ZN(n6098) );
  INV_X1 U3069 ( .A(n6096), .ZN(n6099) );
  INV_X1 U3070 ( .A(n6096), .ZN(n6100) );
  INV_X1 U3071 ( .A(n6096), .ZN(n6101) );
  INV_X1 U3072 ( .A(n6096), .ZN(n6102) );
  INV_X1 U3073 ( .A(n6096), .ZN(n6103) );
  INV_X1 U3074 ( .A(n6105), .ZN(n6106) );
  INV_X1 U3075 ( .A(n6104), .ZN(n6107) );
  INV_X1 U3076 ( .A(n6104), .ZN(n6108) );
  INV_X1 U3077 ( .A(n6104), .ZN(n6109) );
  INV_X1 U3078 ( .A(n6105), .ZN(n6110) );
  INV_X1 U3079 ( .A(n6105), .ZN(n6111) );
  INV_X1 U3080 ( .A(n6116), .ZN(n6117) );
  INV_X1 U3081 ( .A(n6116), .ZN(n6118) );
  INV_X1 U3082 ( .A(n6116), .ZN(n6119) );
  INV_X1 U3083 ( .A(n6116), .ZN(n6120) );
  INV_X1 U3084 ( .A(n6116), .ZN(n6121) );
  INV_X1 U3085 ( .A(n6116), .ZN(n6122) );
  INV_X1 U3086 ( .A(n6116), .ZN(n6123) );
  INV_X1 U3087 ( .A(n6124), .ZN(n6126) );
  INV_X1 U3088 ( .A(n6124), .ZN(n6127) );
  INV_X1 U3089 ( .A(n6125), .ZN(n6128) );
  INV_X1 U3090 ( .A(n6125), .ZN(n6129) );
  INV_X1 U3091 ( .A(n6125), .ZN(n6130) );
  INV_X1 U3092 ( .A(n6124), .ZN(n6131) );
  INV_X1 U3093 ( .A(n2410), .ZN(n6132) );
  INV_X1 U3094 ( .A(n6132), .ZN(n6133) );
  INV_X1 U3095 ( .A(n6132), .ZN(n6134) );
  INV_X1 U3096 ( .A(n6132), .ZN(n6135) );
  INV_X1 U3097 ( .A(n6132), .ZN(n6136) );
  INV_X1 U3098 ( .A(n6132), .ZN(n6137) );
  INV_X1 U3099 ( .A(n6132), .ZN(n6138) );
  INV_X1 U3100 ( .A(n6132), .ZN(n6139) );
  INV_X1 U3101 ( .A(n2412), .ZN(n6140) );
  INV_X1 U3102 ( .A(n6140), .ZN(n6141) );
  INV_X1 U3103 ( .A(n6140), .ZN(n6142) );
  INV_X1 U3104 ( .A(n6140), .ZN(n6143) );
  INV_X1 U3105 ( .A(n6140), .ZN(n6144) );
  INV_X1 U3106 ( .A(n6140), .ZN(n6145) );
  INV_X1 U3107 ( .A(n6140), .ZN(n6146) );
  INV_X1 U3108 ( .A(n6140), .ZN(n6147) );
  INV_X1 U3109 ( .A(n6148), .ZN(n6149) );
  INV_X1 U3110 ( .A(n6148), .ZN(n6150) );
  INV_X1 U3111 ( .A(n6148), .ZN(n6151) );
  INV_X1 U3112 ( .A(n6148), .ZN(n6152) );
  INV_X1 U3113 ( .A(n6148), .ZN(n6153) );
  INV_X1 U3114 ( .A(n6148), .ZN(n6154) );
  INV_X1 U3115 ( .A(n6148), .ZN(n6155) );
  INV_X1 U3116 ( .A(n6156), .ZN(n6158) );
  INV_X1 U3117 ( .A(n6156), .ZN(n6159) );
  INV_X1 U3118 ( .A(n6157), .ZN(n6160) );
  INV_X1 U3119 ( .A(n6157), .ZN(n6161) );
  INV_X1 U3120 ( .A(n6156), .ZN(n6162) );
  INV_X1 U3121 ( .A(n6157), .ZN(n6163) );
  INV_X1 U3122 ( .A(n2403), .ZN(n6164) );
  INV_X1 U3123 ( .A(n6164), .ZN(n6165) );
  INV_X1 U3124 ( .A(n6164), .ZN(n6166) );
  INV_X1 U3125 ( .A(n6164), .ZN(n6167) );
  INV_X1 U3126 ( .A(n6164), .ZN(n6168) );
  INV_X1 U3127 ( .A(n6164), .ZN(n6169) );
  INV_X1 U3128 ( .A(n6164), .ZN(n6170) );
  INV_X1 U3129 ( .A(n6164), .ZN(n6171) );
  INV_X1 U3130 ( .A(n2405), .ZN(n6172) );
  INV_X1 U3131 ( .A(n6172), .ZN(n6173) );
  INV_X1 U3132 ( .A(n6172), .ZN(n6174) );
  INV_X1 U3133 ( .A(n6172), .ZN(n6175) );
  INV_X1 U3134 ( .A(n6172), .ZN(n6176) );
  INV_X1 U3135 ( .A(n6172), .ZN(n6177) );
  INV_X1 U3136 ( .A(n6172), .ZN(n6178) );
  INV_X1 U3137 ( .A(n6172), .ZN(n6179) );
  INV_X1 U3138 ( .A(n6180), .ZN(n6181) );
  INV_X1 U3139 ( .A(n6180), .ZN(n6182) );
  INV_X1 U3140 ( .A(n6180), .ZN(n6183) );
  INV_X1 U3141 ( .A(n6180), .ZN(n6184) );
  INV_X1 U3142 ( .A(n6180), .ZN(n6185) );
  INV_X1 U3143 ( .A(n6180), .ZN(n6186) );
  INV_X1 U3144 ( .A(n6180), .ZN(n6187) );
  INV_X1 U3145 ( .A(n6188), .ZN(n6190) );
  INV_X1 U3146 ( .A(n6188), .ZN(n6191) );
  INV_X1 U3147 ( .A(n6189), .ZN(n6192) );
  INV_X1 U3148 ( .A(n6189), .ZN(n6193) );
  INV_X1 U3149 ( .A(n6188), .ZN(n6194) );
  INV_X1 U3150 ( .A(n6189), .ZN(n6195) );
  INV_X1 U3151 ( .A(n2396), .ZN(n6196) );
  INV_X1 U3152 ( .A(n6196), .ZN(n6197) );
  INV_X1 U3153 ( .A(n6196), .ZN(n6198) );
  INV_X1 U3154 ( .A(n6196), .ZN(n6199) );
  INV_X1 U3155 ( .A(n6196), .ZN(n6200) );
  INV_X1 U3156 ( .A(n6196), .ZN(n6201) );
  INV_X1 U3157 ( .A(n6196), .ZN(n6202) );
  INV_X1 U3158 ( .A(n6196), .ZN(n6203) );
  INV_X1 U3159 ( .A(n2398), .ZN(n6204) );
  INV_X1 U3160 ( .A(n6204), .ZN(n6205) );
  INV_X1 U3161 ( .A(n6204), .ZN(n6206) );
  INV_X1 U3162 ( .A(n6204), .ZN(n6207) );
  INV_X1 U3163 ( .A(n6204), .ZN(n6208) );
  INV_X1 U3164 ( .A(n6204), .ZN(n6209) );
  INV_X1 U3165 ( .A(n6204), .ZN(n6210) );
  INV_X1 U3166 ( .A(n6204), .ZN(n6211) );
  INV_X1 U3167 ( .A(n6212), .ZN(n6213) );
  INV_X1 U3168 ( .A(n6212), .ZN(n6214) );
  INV_X1 U3169 ( .A(n6212), .ZN(n6215) );
  INV_X1 U3170 ( .A(n6212), .ZN(n6216) );
  INV_X1 U3171 ( .A(n6212), .ZN(n6217) );
  INV_X1 U3172 ( .A(n6212), .ZN(n6218) );
  INV_X1 U3173 ( .A(n6212), .ZN(n6219) );
  INV_X1 U3174 ( .A(n6220), .ZN(n6222) );
  INV_X1 U3175 ( .A(n6220), .ZN(n6223) );
  INV_X1 U3176 ( .A(n6221), .ZN(n6224) );
  INV_X1 U3177 ( .A(n6221), .ZN(n6225) );
  INV_X1 U3178 ( .A(n6220), .ZN(n6226) );
  INV_X1 U3179 ( .A(n6221), .ZN(n6227) );
  INV_X1 U3180 ( .A(n2389), .ZN(n6228) );
  INV_X1 U3181 ( .A(n6228), .ZN(n6229) );
  INV_X1 U3182 ( .A(n6228), .ZN(n6230) );
  INV_X1 U3183 ( .A(n6228), .ZN(n6231) );
  INV_X1 U3184 ( .A(n6228), .ZN(n6232) );
  INV_X1 U3185 ( .A(n6228), .ZN(n6233) );
  INV_X1 U3186 ( .A(n6228), .ZN(n6234) );
  INV_X1 U3187 ( .A(n6228), .ZN(n6235) );
  INV_X1 U3188 ( .A(n2391), .ZN(n6236) );
  INV_X1 U3189 ( .A(n6236), .ZN(n6237) );
  INV_X1 U3190 ( .A(n6236), .ZN(n6238) );
  INV_X1 U3191 ( .A(n6236), .ZN(n6239) );
  INV_X1 U3192 ( .A(n6236), .ZN(n6240) );
  INV_X1 U3193 ( .A(n6236), .ZN(n6241) );
  INV_X1 U3194 ( .A(n6236), .ZN(n6242) );
  INV_X1 U3195 ( .A(n6236), .ZN(n6243) );
  INV_X1 U3196 ( .A(n6244), .ZN(n6246) );
  INV_X1 U3197 ( .A(n6244), .ZN(n6247) );
  INV_X1 U3198 ( .A(n6245), .ZN(n6248) );
  INV_X1 U3199 ( .A(n6245), .ZN(n6249) );
  INV_X1 U3200 ( .A(n6245), .ZN(n6250) );
  INV_X1 U3201 ( .A(n6244), .ZN(n6251) );
  INV_X1 U3202 ( .A(n6252), .ZN(n6253) );
  INV_X1 U3203 ( .A(n6252), .ZN(n6254) );
  INV_X1 U3204 ( .A(n6252), .ZN(n6255) );
  INV_X1 U3205 ( .A(n6252), .ZN(n6256) );
  INV_X1 U3206 ( .A(n6252), .ZN(n6257) );
  INV_X1 U3207 ( .A(n6252), .ZN(n6258) );
  INV_X1 U3208 ( .A(n6252), .ZN(n6259) );
  INV_X1 U3209 ( .A(n2378), .ZN(n6260) );
  INV_X1 U3210 ( .A(n6260), .ZN(n6261) );
  INV_X1 U3211 ( .A(n6260), .ZN(n6262) );
  INV_X1 U3212 ( .A(n6260), .ZN(n6263) );
  INV_X1 U3213 ( .A(n6260), .ZN(n6264) );
  INV_X1 U3214 ( .A(n6260), .ZN(n6265) );
  INV_X1 U3215 ( .A(n6260), .ZN(n6266) );
  INV_X1 U3216 ( .A(n6260), .ZN(n6267) );
  INV_X1 U3217 ( .A(n2380), .ZN(n6268) );
  INV_X1 U3218 ( .A(n6268), .ZN(n6269) );
  INV_X1 U3219 ( .A(n6268), .ZN(n6270) );
  INV_X1 U3220 ( .A(n6268), .ZN(n6271) );
  INV_X1 U3221 ( .A(n6268), .ZN(n6272) );
  INV_X1 U3222 ( .A(n6268), .ZN(n6273) );
  INV_X1 U3223 ( .A(n6268), .ZN(n6274) );
  INV_X1 U3224 ( .A(n6268), .ZN(n6275) );
  INV_X1 U3225 ( .A(n6276), .ZN(n6278) );
  INV_X1 U3226 ( .A(n6276), .ZN(n6279) );
  INV_X1 U3227 ( .A(n6277), .ZN(n6280) );
  INV_X1 U3228 ( .A(n6277), .ZN(n6281) );
  INV_X1 U3229 ( .A(n6277), .ZN(n6282) );
  INV_X1 U3230 ( .A(n6276), .ZN(n6283) );
  INV_X1 U3231 ( .A(n6284), .ZN(n6285) );
  INV_X1 U3232 ( .A(n6284), .ZN(n6286) );
  INV_X1 U3233 ( .A(n6284), .ZN(n6287) );
  INV_X1 U3234 ( .A(n6284), .ZN(n6288) );
  INV_X1 U3235 ( .A(n6284), .ZN(n6289) );
  INV_X1 U3236 ( .A(n6284), .ZN(n6290) );
  INV_X1 U3237 ( .A(n6284), .ZN(n6291) );
  INV_X1 U3238 ( .A(n2371), .ZN(n6292) );
  INV_X1 U3239 ( .A(n6292), .ZN(n6293) );
  INV_X1 U3240 ( .A(n6292), .ZN(n6294) );
  INV_X1 U3241 ( .A(n6292), .ZN(n6295) );
  INV_X1 U3242 ( .A(n6292), .ZN(n6296) );
  INV_X1 U3243 ( .A(n6292), .ZN(n6297) );
  INV_X1 U3244 ( .A(n6292), .ZN(n6298) );
  INV_X1 U3245 ( .A(n6292), .ZN(n6299) );
  INV_X1 U3246 ( .A(n2373), .ZN(n6300) );
  INV_X1 U3247 ( .A(n6300), .ZN(n6301) );
  INV_X1 U3248 ( .A(n6300), .ZN(n6302) );
  INV_X1 U3249 ( .A(n6300), .ZN(n6303) );
  INV_X1 U3250 ( .A(n6300), .ZN(n6304) );
  INV_X1 U3251 ( .A(n6300), .ZN(n6305) );
  INV_X1 U3252 ( .A(n6300), .ZN(n6306) );
  INV_X1 U3253 ( .A(n6300), .ZN(n6307) );
  INV_X1 U3254 ( .A(n6308), .ZN(n6309) );
  INV_X1 U3255 ( .A(n6308), .ZN(n6310) );
  INV_X1 U3256 ( .A(n6308), .ZN(n6311) );
  INV_X1 U3257 ( .A(n6308), .ZN(n6312) );
  INV_X1 U3258 ( .A(n6308), .ZN(n6313) );
  INV_X1 U3259 ( .A(n6308), .ZN(n6314) );
  INV_X1 U3260 ( .A(n6308), .ZN(n6315) );
  INV_X1 U3261 ( .A(n6316), .ZN(n6318) );
  INV_X1 U3262 ( .A(n6316), .ZN(n6319) );
  INV_X1 U3263 ( .A(n6317), .ZN(n6320) );
  INV_X1 U3264 ( .A(n6317), .ZN(n6321) );
  INV_X1 U3265 ( .A(n6316), .ZN(n6322) );
  INV_X1 U3266 ( .A(n6317), .ZN(n6323) );
  INV_X1 U3267 ( .A(n6328), .ZN(n6329) );
  INV_X1 U3268 ( .A(n6328), .ZN(n6330) );
  INV_X1 U3269 ( .A(n6328), .ZN(n6331) );
  INV_X1 U3270 ( .A(n6328), .ZN(n6332) );
  INV_X1 U3271 ( .A(n6328), .ZN(n6333) );
  INV_X1 U3272 ( .A(n6328), .ZN(n6334) );
  INV_X1 U3273 ( .A(n6328), .ZN(n6335) );
  INV_X1 U3274 ( .A(n6336), .ZN(n6338) );
  INV_X1 U3275 ( .A(n6336), .ZN(n6339) );
  INV_X1 U3276 ( .A(n6337), .ZN(n6340) );
  INV_X1 U3277 ( .A(n6337), .ZN(n6341) );
  INV_X1 U3278 ( .A(n6336), .ZN(n6342) );
  INV_X1 U3279 ( .A(n6337), .ZN(n6343) );
  INV_X1 U3280 ( .A(n6736), .ZN(n6734) );
  INV_X1 U3281 ( .A(n6736), .ZN(n6735) );
endmodule


module FETCH_UNIT_NB32_LS5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , n1;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X1 U2 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  XOR2_X1 U5 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  XOR2_X1 U7 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  XOR2_X1 U9 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  XOR2_X1 U11 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  XOR2_X1 U13 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  XOR2_X1 U15 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  XOR2_X1 U17 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  XOR2_X1 U19 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  XOR2_X1 U21 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X1 U25 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  XOR2_X1 U27 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  XOR2_X1 U29 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  XOR2_X1 U31 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  XOR2_X1 U33 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  XOR2_X1 U35 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  XOR2_X1 U37 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  XOR2_X1 U39 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  XOR2_X1 U41 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  XOR2_X1 U43 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  XOR2_X1 U45 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  XOR2_X1 U47 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  XOR2_X1 U49 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  XOR2_X1 U51 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  XOR2_X1 U53 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U55 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  XOR2_X1 U57 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  XNOR2_X1 U1 ( .A(A[31]), .B(n1), .ZN(SUM[31]) );
  NAND2_X1 U3 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n1) );
  INV_X1 U4 ( .A(\carry[3] ), .ZN(SUM[2]) );
  AND2_X1 U6 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  AND2_X1 U8 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  AND2_X1 U10 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  AND2_X1 U12 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  AND2_X1 U14 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  AND2_X1 U16 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  AND2_X1 U18 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  AND2_X1 U20 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  AND2_X1 U22 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  AND2_X1 U24 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  AND2_X1 U26 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  AND2_X1 U28 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  AND2_X1 U30 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  AND2_X1 U32 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  AND2_X1 U34 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  AND2_X1 U36 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U38 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U40 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  AND2_X1 U42 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  AND2_X1 U44 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  AND2_X1 U46 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  AND2_X1 U48 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  AND2_X1 U50 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  AND2_X1 U52 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  AND2_X1 U54 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  AND2_X1 U56 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  AND2_X1 U58 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
endmodule


module MUX21_generic_NB32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77;

  INV_X1 U1 ( .A(n76), .ZN(n67) );
  BUF_X1 U2 ( .A(n77), .Z(n73) );
  BUF_X1 U3 ( .A(n77), .Z(n68) );
  BUF_X1 U4 ( .A(n77), .Z(n76) );
  BUF_X1 U5 ( .A(n73), .Z(n74) );
  BUF_X1 U6 ( .A(n77), .Z(n69) );
  BUF_X1 U7 ( .A(n70), .Z(n75) );
  BUF_X1 U8 ( .A(n77), .Z(n72) );
  BUF_X1 U9 ( .A(n77), .Z(n71) );
  BUF_X1 U10 ( .A(n77), .Z(n70) );
  INV_X1 U11 ( .A(n53), .ZN(Y[21]) );
  INV_X1 U12 ( .A(n34), .ZN(Y[9]) );
  INV_X1 U13 ( .A(n60), .ZN(Y[15]) );
  INV_X1 U14 ( .A(n47), .ZN(Y[27]) );
  INV_X1 U15 ( .A(n42), .ZN(Y[31]) );
  INV_X1 U16 ( .A(n64), .ZN(Y[11]) );
  INV_X1 U17 ( .A(n65), .ZN(Y[10]) );
  INV_X1 U18 ( .A(n41), .ZN(Y[3]) );
  INV_X1 U19 ( .A(n40), .ZN(Y[4]) );
  INV_X1 U20 ( .A(n38), .ZN(Y[6]) );
  INV_X1 U21 ( .A(n37), .ZN(Y[7]) );
  INV_X1 U22 ( .A(n61), .ZN(Y[14]) );
  INV_X1 U23 ( .A(n57), .ZN(Y[18]) );
  INV_X1 U24 ( .A(n52), .ZN(Y[22]) );
  INV_X1 U25 ( .A(n48), .ZN(Y[26]) );
  INV_X1 U26 ( .A(n62), .ZN(Y[13]) );
  INV_X1 U27 ( .A(n44), .ZN(Y[2]) );
  INV_X1 U28 ( .A(n39), .ZN(Y[5]) );
  INV_X1 U29 ( .A(n56), .ZN(Y[19]) );
  INV_X1 U30 ( .A(n54), .ZN(Y[20]) );
  INV_X1 U31 ( .A(n51), .ZN(Y[23]) );
  INV_X1 U32 ( .A(n50), .ZN(Y[24]) );
  INV_X1 U33 ( .A(n49), .ZN(Y[25]) );
  INV_X1 U34 ( .A(n46), .ZN(Y[28]) );
  INV_X1 U35 ( .A(n45), .ZN(Y[29]) );
  INV_X1 U36 ( .A(n63), .ZN(Y[12]) );
  INV_X1 U37 ( .A(n59), .ZN(Y[16]) );
  INV_X1 U38 ( .A(n58), .ZN(Y[17]) );
  INV_X1 U39 ( .A(n36), .ZN(Y[8]) );
  AOI22_X1 U40 ( .A1(SEL), .A2(A[9]), .B1(B[9]), .B2(n68), .ZN(n34) );
  AOI22_X1 U41 ( .A1(A[10]), .A2(n67), .B1(B[10]), .B2(n75), .ZN(n65) );
  AOI22_X1 U42 ( .A1(A[11]), .A2(n67), .B1(B[11]), .B2(n75), .ZN(n64) );
  AOI22_X1 U43 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(n69), .ZN(n41) );
  AOI22_X1 U44 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(n69), .ZN(n40) );
  AOI22_X1 U45 ( .A1(A[6]), .A2(SEL), .B1(B[6]), .B2(n68), .ZN(n38) );
  AOI22_X1 U46 ( .A1(A[7]), .A2(SEL), .B1(B[7]), .B2(n68), .ZN(n37) );
  AOI22_X1 U47 ( .A1(A[14]), .A2(n67), .B1(B[14]), .B2(n74), .ZN(n61) );
  AOI22_X1 U48 ( .A1(A[19]), .A2(n67), .B1(B[19]), .B2(n73), .ZN(n56) );
  AOI22_X1 U49 ( .A1(A[5]), .A2(SEL), .B1(B[5]), .B2(n69), .ZN(n39) );
  AOI22_X1 U50 ( .A1(A[8]), .A2(n67), .B1(B[8]), .B2(n68), .ZN(n36) );
  AOI22_X1 U51 ( .A1(A[15]), .A2(n67), .B1(B[15]), .B2(n74), .ZN(n60) );
  AOI22_X1 U52 ( .A1(A[16]), .A2(n67), .B1(B[16]), .B2(n74), .ZN(n59) );
  AOI22_X1 U53 ( .A1(A[17]), .A2(n67), .B1(B[17]), .B2(n73), .ZN(n58) );
  AOI22_X1 U54 ( .A1(A[18]), .A2(n67), .B1(B[18]), .B2(n73), .ZN(n57) );
  AOI22_X1 U55 ( .A1(A[22]), .A2(SEL), .B1(B[22]), .B2(n72), .ZN(n52) );
  AOI22_X1 U56 ( .A1(A[23]), .A2(SEL), .B1(B[23]), .B2(n72), .ZN(n51) );
  AOI22_X1 U57 ( .A1(A[27]), .A2(SEL), .B1(B[27]), .B2(n71), .ZN(n47) );
  AOI22_X1 U58 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n70), .ZN(n44) );
  INV_X1 U59 ( .A(SEL), .ZN(n77) );
  INV_X1 U60 ( .A(n66), .ZN(Y[0]) );
  INV_X1 U61 ( .A(n55), .ZN(Y[1]) );
  AOI22_X1 U62 ( .A1(A[0]), .A2(n67), .B1(B[0]), .B2(n75), .ZN(n66) );
  AOI22_X1 U63 ( .A1(A[1]), .A2(n67), .B1(B[1]), .B2(n73), .ZN(n55) );
  AOI22_X1 U64 ( .A1(A[12]), .A2(n67), .B1(B[12]), .B2(n75), .ZN(n63) );
  AOI22_X1 U65 ( .A1(A[30]), .A2(SEL), .B1(B[30]), .B2(n70), .ZN(n43) );
  INV_X1 U66 ( .A(n43), .ZN(Y[30]) );
  AOI22_X1 U67 ( .A1(A[28]), .A2(SEL), .B1(B[28]), .B2(n70), .ZN(n46) );
  AOI22_X1 U68 ( .A1(A[25]), .A2(SEL), .B1(B[25]), .B2(n71), .ZN(n49) );
  AOI22_X1 U69 ( .A1(A[20]), .A2(SEL), .B1(B[20]), .B2(n72), .ZN(n54) );
  AOI22_X1 U70 ( .A1(A[26]), .A2(SEL), .B1(B[26]), .B2(n71), .ZN(n48) );
  AOI22_X1 U71 ( .A1(A[31]), .A2(n67), .B1(B[31]), .B2(n69), .ZN(n42) );
  AOI22_X1 U72 ( .A1(A[24]), .A2(n67), .B1(B[24]), .B2(n71), .ZN(n50) );
  AOI22_X1 U73 ( .A1(A[13]), .A2(n67), .B1(B[13]), .B2(n74), .ZN(n62) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n67), .B1(B[29]), .B2(n70), .ZN(n45) );
  AOI22_X1 U75 ( .A1(A[21]), .A2(SEL), .B1(B[21]), .B2(n72), .ZN(n53) );
endmodule


module FD_NB32_5 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n35, n68, n69, n70;
  assign n35 = RESET;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n70), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n70), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n70), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n70), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n70), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n70), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n70), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n70), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n68), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n68), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n68), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n68), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n68), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n68), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n68), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n68), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n68), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n68), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n68), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n68), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n69), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n69), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n69), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n69), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n69), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n69), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n69), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n69), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n69), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n69), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n69), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n69), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n35), .Z(n69) );
  BUF_X1 U4 ( .A(n35), .Z(n68) );
  BUF_X1 U5 ( .A(n35), .Z(n70) );
endmodule


module MUX21_generic_NB32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n39, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82;

  CLKBUF_X1 U1 ( .A(n82), .Z(n74) );
  BUF_X1 U2 ( .A(n82), .Z(n81) );
  BUF_X1 U3 ( .A(n82), .Z(n73) );
  BUF_X1 U4 ( .A(n79), .Z(n77) );
  BUF_X1 U5 ( .A(n79), .Z(n76) );
  BUF_X1 U6 ( .A(SEL), .Z(n70) );
  INV_X1 U7 ( .A(B[5]), .ZN(n69) );
  INV_X1 U8 ( .A(A[5]), .ZN(n68) );
  INV_X1 U9 ( .A(n65), .ZN(Y[10]) );
  INV_X1 U10 ( .A(n64), .ZN(Y[11]) );
  INV_X1 U11 ( .A(n38), .ZN(Y[6]) );
  INV_X1 U12 ( .A(n40), .ZN(Y[4]) );
  INV_X1 U13 ( .A(n62), .ZN(Y[13]) );
  INV_X1 U14 ( .A(n61), .ZN(Y[14]) );
  INV_X1 U15 ( .A(n63), .ZN(Y[12]) );
  INV_X1 U16 ( .A(n43), .ZN(Y[30]) );
  INV_X1 U17 ( .A(n45), .ZN(Y[29]) );
  INV_X1 U18 ( .A(n42), .ZN(Y[31]) );
  INV_X1 U19 ( .A(n47), .ZN(Y[27]) );
  INV_X1 U20 ( .A(n46), .ZN(Y[28]) );
  INV_X1 U21 ( .A(n60), .ZN(Y[15]) );
  INV_X1 U22 ( .A(n59), .ZN(Y[16]) );
  INV_X1 U23 ( .A(n58), .ZN(Y[17]) );
  INV_X1 U24 ( .A(n57), .ZN(Y[18]) );
  INV_X1 U25 ( .A(n56), .ZN(Y[19]) );
  INV_X1 U26 ( .A(n54), .ZN(Y[20]) );
  INV_X1 U27 ( .A(n53), .ZN(Y[21]) );
  INV_X1 U28 ( .A(n52), .ZN(Y[22]) );
  INV_X1 U29 ( .A(n51), .ZN(Y[23]) );
  INV_X1 U30 ( .A(n50), .ZN(Y[24]) );
  INV_X1 U31 ( .A(n49), .ZN(Y[25]) );
  INV_X1 U32 ( .A(n48), .ZN(Y[26]) );
  CLKBUF_X1 U33 ( .A(n74), .Z(n79) );
  CLKBUF_X1 U34 ( .A(n82), .Z(n80) );
  INV_X1 U35 ( .A(n41), .ZN(Y[3]) );
  INV_X1 U36 ( .A(n82), .ZN(n39) );
  INV_X1 U37 ( .A(n34), .ZN(Y[9]) );
  INV_X1 U38 ( .A(n37), .ZN(Y[7]) );
  INV_X1 U39 ( .A(n66), .ZN(Y[0]) );
  INV_X1 U40 ( .A(n36), .ZN(Y[8]) );
  OAI22_X1 U41 ( .A1(n68), .A2(n74), .B1(n69), .B2(n72), .ZN(Y[5]) );
  INV_X2 U42 ( .A(n81), .ZN(n72) );
  CLKBUF_X1 U43 ( .A(n82), .Z(n75) );
  INV_X1 U44 ( .A(n70), .ZN(n82) );
  AOI22_X1 U45 ( .A1(A[20]), .A2(n71), .B1(B[20]), .B2(n77), .ZN(n54) );
  AOI22_X1 U46 ( .A1(A[25]), .A2(n72), .B1(B[25]), .B2(n76), .ZN(n49) );
  AOI22_X1 U47 ( .A1(A[24]), .A2(n71), .B1(B[24]), .B2(n76), .ZN(n50) );
  AOI22_X1 U48 ( .A1(A[21]), .A2(n71), .B1(B[21]), .B2(n77), .ZN(n53) );
  AOI22_X1 U49 ( .A1(A[22]), .A2(n71), .B1(B[22]), .B2(n77), .ZN(n52) );
  AOI22_X1 U50 ( .A1(A[26]), .A2(n72), .B1(B[26]), .B2(n76), .ZN(n48) );
  AOI22_X1 U51 ( .A1(A[23]), .A2(n71), .B1(B[23]), .B2(n77), .ZN(n51) );
  AOI22_X1 U52 ( .A1(A[28]), .A2(n72), .B1(B[28]), .B2(n75), .ZN(n46) );
  AOI22_X1 U53 ( .A1(A[27]), .A2(n71), .B1(B[27]), .B2(n76), .ZN(n47) );
  AOI22_X1 U54 ( .A1(A[29]), .A2(n71), .B1(B[29]), .B2(n75), .ZN(n45) );
  AOI22_X1 U55 ( .A1(A[30]), .A2(n72), .B1(B[30]), .B2(n75), .ZN(n43) );
  INV_X1 U56 ( .A(n44), .ZN(Y[2]) );
  AOI22_X1 U57 ( .A1(A[2]), .A2(n39), .B1(B[2]), .B2(n75), .ZN(n44) );
  INV_X1 U58 ( .A(n55), .ZN(Y[1]) );
  BUF_X1 U59 ( .A(n73), .Z(n78) );
  INV_X2 U60 ( .A(n81), .ZN(n71) );
  AOI22_X1 U61 ( .A1(A[17]), .A2(n72), .B1(B[17]), .B2(n78), .ZN(n58) );
  AOI22_X1 U62 ( .A1(A[18]), .A2(n71), .B1(B[18]), .B2(n78), .ZN(n57) );
  AOI22_X1 U63 ( .A1(A[16]), .A2(n72), .B1(B[16]), .B2(n79), .ZN(n59) );
  AOI22_X1 U64 ( .A1(A[19]), .A2(n72), .B1(B[19]), .B2(n78), .ZN(n56) );
  AOI22_X1 U65 ( .A1(A[14]), .A2(n71), .B1(B[14]), .B2(n79), .ZN(n61) );
  AOI22_X1 U66 ( .A1(A[12]), .A2(n71), .B1(B[12]), .B2(n80), .ZN(n63) );
  AOI22_X1 U67 ( .A1(A[13]), .A2(n71), .B1(B[13]), .B2(n79), .ZN(n62) );
  AOI22_X1 U68 ( .A1(A[15]), .A2(n71), .B1(B[15]), .B2(n79), .ZN(n60) );
  AOI22_X1 U69 ( .A1(A[11]), .A2(n71), .B1(B[11]), .B2(n80), .ZN(n64) );
  AOI22_X1 U70 ( .A1(A[10]), .A2(n72), .B1(B[10]), .B2(n80), .ZN(n65) );
  AOI22_X1 U71 ( .A1(A[0]), .A2(n39), .B1(B[0]), .B2(n80), .ZN(n66) );
  AOI22_X1 U72 ( .A1(A[1]), .A2(n39), .B1(B[1]), .B2(n78), .ZN(n55) );
  AOI22_X1 U73 ( .A1(A[31]), .A2(n72), .B1(B[31]), .B2(n74), .ZN(n42) );
  AOI22_X1 U74 ( .A1(A[8]), .A2(n71), .B1(B[8]), .B2(n73), .ZN(n36) );
  AOI22_X1 U75 ( .A1(A[3]), .A2(n72), .B1(B[3]), .B2(n74), .ZN(n41) );
  AOI22_X1 U76 ( .A1(A[7]), .A2(n72), .B1(B[7]), .B2(n73), .ZN(n37) );
  AOI22_X1 U77 ( .A1(n39), .A2(A[9]), .B1(B[9]), .B2(n73), .ZN(n34) );
  AOI22_X1 U78 ( .A1(A[6]), .A2(n39), .B1(B[6]), .B2(n73), .ZN(n38) );
  AOI22_X1 U79 ( .A1(A[4]), .A2(n39), .B1(B[4]), .B2(n74), .ZN(n40) );
endmodule


module FD_NB32_0 ( CK, RESET, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n35, n36, n37, n38;
  assign n35 = RESET;

  DFFR_X1 \TMP_Q_reg[31]  ( .D(D[31]), .CK(CK), .RN(n38), .Q(Q[31]) );
  DFFR_X1 \TMP_Q_reg[30]  ( .D(D[30]), .CK(CK), .RN(n38), .Q(Q[30]) );
  DFFR_X1 \TMP_Q_reg[29]  ( .D(D[29]), .CK(CK), .RN(n38), .Q(Q[29]) );
  DFFR_X1 \TMP_Q_reg[28]  ( .D(D[28]), .CK(CK), .RN(n38), .Q(Q[28]) );
  DFFR_X1 \TMP_Q_reg[27]  ( .D(D[27]), .CK(CK), .RN(n38), .Q(Q[27]) );
  DFFR_X1 \TMP_Q_reg[26]  ( .D(D[26]), .CK(CK), .RN(n38), .Q(Q[26]) );
  DFFR_X1 \TMP_Q_reg[25]  ( .D(D[25]), .CK(CK), .RN(n38), .Q(Q[25]) );
  DFFR_X1 \TMP_Q_reg[24]  ( .D(D[24]), .CK(CK), .RN(n38), .Q(Q[24]) );
  DFFR_X1 \TMP_Q_reg[23]  ( .D(D[23]), .CK(CK), .RN(n36), .Q(Q[23]) );
  DFFR_X1 \TMP_Q_reg[22]  ( .D(D[22]), .CK(CK), .RN(n36), .Q(Q[22]) );
  DFFR_X1 \TMP_Q_reg[21]  ( .D(D[21]), .CK(CK), .RN(n36), .Q(Q[21]) );
  DFFR_X1 \TMP_Q_reg[20]  ( .D(D[20]), .CK(CK), .RN(n36), .Q(Q[20]) );
  DFFR_X1 \TMP_Q_reg[19]  ( .D(D[19]), .CK(CK), .RN(n36), .Q(Q[19]) );
  DFFR_X1 \TMP_Q_reg[18]  ( .D(D[18]), .CK(CK), .RN(n36), .Q(Q[18]) );
  DFFR_X1 \TMP_Q_reg[17]  ( .D(D[17]), .CK(CK), .RN(n36), .Q(Q[17]) );
  DFFR_X1 \TMP_Q_reg[16]  ( .D(D[16]), .CK(CK), .RN(n36), .Q(Q[16]) );
  DFFR_X1 \TMP_Q_reg[15]  ( .D(D[15]), .CK(CK), .RN(n36), .Q(Q[15]) );
  DFFR_X1 \TMP_Q_reg[14]  ( .D(D[14]), .CK(CK), .RN(n36), .Q(Q[14]) );
  DFFR_X1 \TMP_Q_reg[13]  ( .D(D[13]), .CK(CK), .RN(n36), .Q(Q[13]) );
  DFFR_X1 \TMP_Q_reg[12]  ( .D(D[12]), .CK(CK), .RN(n36), .Q(Q[12]) );
  DFFR_X1 \TMP_Q_reg[11]  ( .D(D[11]), .CK(CK), .RN(n37), .Q(Q[11]) );
  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(n37), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(n37), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(n37), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(n37), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(n37), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(n37), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(n37), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(n37), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(n37), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(n37), .Q(Q[0]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(n37), .Q(Q[1]) );
  BUF_X1 U3 ( .A(n35), .Z(n37) );
  BUF_X1 U4 ( .A(n35), .Z(n36) );
  BUF_X1 U5 ( .A(n35), .Z(n38) );
endmodule


module BP_NB32_BP_LEN4 ( CLK, RST, EX_PC, CURR_PC, NEXT_PC, NEW_PC, INST, 
        MISS_HIT, PRED );
  input [31:0] EX_PC;
  input [31:0] CURR_PC;
  input [31:0] NEXT_PC;
  input [31:0] NEW_PC;
  input [31:0] INST;
  output [1:0] MISS_HIT;
  output [31:0] PRED;
  input CLK, RST;
  wire   INST_31, INST_30, INST_29, INST_28, INST_27, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, \PRED_HISTORY[0][32] ,
         \PRED_HISTORY[0][31] , \PRED_HISTORY[0][30] , \PRED_HISTORY[0][29] ,
         \PRED_HISTORY[0][28] , \PRED_HISTORY[0][27] , \PRED_HISTORY[0][26] ,
         \PRED_HISTORY[0][25] , \PRED_HISTORY[0][24] , \PRED_HISTORY[0][23] ,
         \PRED_HISTORY[0][22] , \PRED_HISTORY[0][21] , \PRED_HISTORY[0][20] ,
         \PRED_HISTORY[0][19] , \PRED_HISTORY[0][18] , \PRED_HISTORY[0][17] ,
         \PRED_HISTORY[0][16] , \PRED_HISTORY[0][15] , \PRED_HISTORY[0][14] ,
         \PRED_HISTORY[0][13] , \PRED_HISTORY[0][12] , \PRED_HISTORY[0][11] ,
         \PRED_HISTORY[0][10] , \PRED_HISTORY[0][9] , \PRED_HISTORY[0][8] ,
         \PRED_HISTORY[0][7] , \PRED_HISTORY[0][6] , \PRED_HISTORY[0][5] ,
         \PRED_HISTORY[0][4] , \PRED_HISTORY[0][3] , \PRED_HISTORY[0][2] ,
         \PRED_HISTORY[0][1] , \PRED_HISTORY[0][0] , \PRED_HISTORY[1][31] ,
         \PRED_HISTORY[1][30] , \PRED_HISTORY[1][29] , \PRED_HISTORY[1][28] ,
         \PRED_HISTORY[1][27] , \PRED_HISTORY[1][26] , \PRED_HISTORY[1][25] ,
         \PRED_HISTORY[1][24] , \PRED_HISTORY[1][23] , \PRED_HISTORY[1][22] ,
         \PRED_HISTORY[1][21] , \PRED_HISTORY[1][20] , \PRED_HISTORY[1][19] ,
         \PRED_HISTORY[1][18] , \PRED_HISTORY[1][17] , \PRED_HISTORY[1][16] ,
         \PRED_HISTORY[1][15] , \PRED_HISTORY[1][14] , \PRED_HISTORY[1][13] ,
         \PRED_HISTORY[1][12] , \PRED_HISTORY[1][11] , \PRED_HISTORY[1][10] ,
         \PRED_HISTORY[1][9] , \PRED_HISTORY[1][8] , \PRED_HISTORY[1][7] ,
         \PRED_HISTORY[1][6] , \PRED_HISTORY[1][5] , \PRED_HISTORY[1][4] ,
         \PRED_HISTORY[1][3] , \PRED_HISTORY[1][2] , \PRED_HISTORY[1][1] ,
         \PRED_HISTORY[1][0] , N815, \PC_HISTORY[0][3] , \PC_HISTORY[0][2] ,
         \PC_HISTORY[0][1] , \PC_HISTORY[0][0] , n194, n197, n198, n210, n213,
         n214, n226, n229, n230, n242, n245, n246, n258, n261, n262, n274,
         n277, n278, n290, n293, n294, n306, n309, n310, n322, n325, n326,
         n338, n341, n342, n354, n357, n358, n361, n370, n373, n374, n390,
         n418, n450, n453, n454, n466, n469, n470, n482, n485, n486, n498,
         n501, n502, n514, n517, n518, n530, n533, n534, n546, n549, n550,
         n562, n565, n566, n578, n581, n582, n594, n597, n598, n610, n613,
         n614, n626, n629, n630, n642, n645, n646, n658, n661, n662, n674,
         n677, n678, n690, n699, n700, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n818, n819, n820, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n834, n835,
         n836, n837, n838, n839, n842, n843, n844, n846, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n863, n864, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n958, n959, n960, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n991,
         n992, n994, n995, n996, n997, n998, n999, n1068, n1070, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1360,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1476, n1477, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1571, n1572, n1573,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1604, n1605, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1668, n1669,
         n1670, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1732, n1733,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1763, n1764, n1765, n1766,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1796, n1797, n1798, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1827, n1828, n1829, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1860, n1861, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n3, n4, n5, n6, n7, n9, n42, n43, n44, n52, n55, n56, n58, n59, n61,
         n88, n89, n92, n96, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n1411, n1446, n1475, n1478, n1506, n1538, n1539, n1570, n1795,
         n1799, n1826, n1830, n1831, n1858, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1918, n1940, n1941, n1942, n1943,
         n1958, n1959, n1960, n1961, n2246, n2362, n2048, n2049, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2210, n2211, n2213, n2215,
         n2217, n2219, n2221, n2223, n2225, n2227, n2229, n2231, n2233, n2235,
         n2237, n2239, n2243, n2245, n2248, n2250, n2252, n2254, n2256, n2258,
         n2260, n2262, n2264, n2266, n2268, n2269, n2270, n2271, n2298, n2299,
         n2300, n2332, n2333, n2335, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2448, n2449, n2452, n2453,
         n2454, n2456, n2459, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2473, n2474, n2475, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2499, n2500,
         n2501, n2502, n2504, n2505, n2508, n2509, n2510, n2511, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2654, n2656, n2657, n2658, n2659,
         n2660, n2661, n2663, n2664, n2665, n2667, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2412, n2421, n2447, n2450, n2451, n2455,
         n2457, n2458, n2460, n2472, n2476, n2498, n2503, n2506, n2507, n2512,
         n2513, n2514, n2522, n2535, n2546, n2557, n2568, n2579, n2590, n2601,
         n2612, n2623, n2644, n2653, n2655, n2662, n2666, n2668, n2679, n2690,
         n2701, n2712, n2723, n2734, n2745, n2756, n2767, n2789, n2800, n2811,
         n2822, n2833, n2844, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2968, n2969, n2970, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245;
  wire   [31:0] PRED_TK;
  assign INST_31 = INST[31];
  assign INST_30 = INST[30];
  assign INST_29 = INST[29];
  assign INST_28 = INST[28];
  assign INST_27 = INST[27];
  assign n2246 = RST;

  DFFR_X1 \PRED_HISTORY_reg[0][32]  ( .D(n2362), .CK(CLK), .RN(n3202), .Q(
        \PRED_HISTORY[0][32] ) );
  DFFR_X1 \PC_HISTORY_reg[0][3]  ( .D(CURR_PC[5]), .CK(CLK), .RN(n3203), .Q(
        \PC_HISTORY[0][3] ) );
  DFFR_X1 \PC_HISTORY_reg[0][2]  ( .D(CURR_PC[4]), .CK(CLK), .RN(n3203), .Q(
        \PC_HISTORY[0][2] ) );
  DFFR_X1 \PC_HISTORY_reg[0][1]  ( .D(CURR_PC[3]), .CK(CLK), .RN(n3221), .Q(
        \PC_HISTORY[0][1] ) );
  DFFR_X1 \PC_HISTORY_reg[0][0]  ( .D(CURR_PC[2]), .CK(CLK), .RN(n3221), .Q(
        \PC_HISTORY[0][0] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][0]  ( .D(PRED[0]), .CK(CLK), .RN(n3221), .Q(
        \PRED_HISTORY[0][0] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][0]  ( .D(\PRED_HISTORY[0][0] ), .CK(CLK), .RN(
        n3221), .Q(\PRED_HISTORY[1][0] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][9]  ( .D(PRED[9]), .CK(CLK), .RN(n3221), .Q(
        \PRED_HISTORY[0][9] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][9]  ( .D(\PRED_HISTORY[0][9] ), .CK(CLK), .RN(
        n3221), .Q(\PRED_HISTORY[1][9] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][8]  ( .D(PRED[8]), .CK(CLK), .RN(n3221), .Q(
        \PRED_HISTORY[0][8] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][8]  ( .D(\PRED_HISTORY[0][8] ), .CK(CLK), .RN(
        n3202), .Q(\PRED_HISTORY[1][8] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][7]  ( .D(PRED[7]), .CK(CLK), .RN(n3202), .Q(
        \PRED_HISTORY[0][7] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][7]  ( .D(\PRED_HISTORY[0][7] ), .CK(CLK), .RN(
        n3202), .Q(\PRED_HISTORY[1][7] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][6]  ( .D(PRED[6]), .CK(CLK), .RN(n3202), .Q(
        \PRED_HISTORY[0][6] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][6]  ( .D(\PRED_HISTORY[0][6] ), .CK(CLK), .RN(
        n3202), .Q(\PRED_HISTORY[1][6] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][5]  ( .D(PRED[5]), .CK(CLK), .RN(n3202), .Q(
        \PRED_HISTORY[0][5] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][5]  ( .D(\PRED_HISTORY[0][5] ), .CK(CLK), .RN(
        n3202), .Q(\PRED_HISTORY[1][5] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][4]  ( .D(PRED[4]), .CK(CLK), .RN(n3201), .Q(
        \PRED_HISTORY[0][4] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][4]  ( .D(\PRED_HISTORY[0][4] ), .CK(CLK), .RN(
        n3202), .Q(\PRED_HISTORY[1][4] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][3]  ( .D(PRED[3]), .CK(CLK), .RN(n3202), .Q(
        \PRED_HISTORY[0][3] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][3]  ( .D(\PRED_HISTORY[0][3] ), .CK(CLK), .RN(
        n3202), .Q(\PRED_HISTORY[1][3] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][31]  ( .D(PRED[31]), .CK(CLK), .RN(n3202), .Q(
        \PRED_HISTORY[0][31] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][31]  ( .D(\PRED_HISTORY[0][31] ), .CK(CLK), 
        .RN(n3222), .Q(\PRED_HISTORY[1][31] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][30]  ( .D(PRED[30]), .CK(CLK), .RN(n3221), .Q(
        \PRED_HISTORY[0][30] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][30]  ( .D(\PRED_HISTORY[0][30] ), .CK(CLK), 
        .RN(n3221), .Q(\PRED_HISTORY[1][30] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][2]  ( .D(PRED[2]), .CK(CLK), .RN(n3222), .Q(
        \PRED_HISTORY[0][2] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][2]  ( .D(\PRED_HISTORY[0][2] ), .CK(CLK), .RN(
        n3222), .Q(\PRED_HISTORY[1][2] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][29]  ( .D(PRED[29]), .CK(CLK), .RN(n3222), .Q(
        \PRED_HISTORY[0][29] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][29]  ( .D(\PRED_HISTORY[0][29] ), .CK(CLK), 
        .RN(n3222), .Q(\PRED_HISTORY[1][29] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][28]  ( .D(PRED[28]), .CK(CLK), .RN(n3222), .Q(
        \PRED_HISTORY[0][28] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][28]  ( .D(\PRED_HISTORY[0][28] ), .CK(CLK), 
        .RN(n3222), .Q(\PRED_HISTORY[1][28] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][27]  ( .D(PRED[27]), .CK(CLK), .RN(n3222), .Q(
        \PRED_HISTORY[0][27] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][27]  ( .D(\PRED_HISTORY[0][27] ), .CK(CLK), 
        .RN(n3222), .Q(\PRED_HISTORY[1][27] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][26]  ( .D(PRED[26]), .CK(CLK), .RN(n3222), .Q(
        \PRED_HISTORY[0][26] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][26]  ( .D(\PRED_HISTORY[0][26] ), .CK(CLK), 
        .RN(n3201), .Q(\PRED_HISTORY[1][26] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][25]  ( .D(PRED[25]), .CK(CLK), .RN(n3201), .Q(
        \PRED_HISTORY[0][25] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][25]  ( .D(\PRED_HISTORY[0][25] ), .CK(CLK), 
        .RN(n3201), .Q(\PRED_HISTORY[1][25] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][24]  ( .D(PRED[24]), .CK(CLK), .RN(n3201), .Q(
        \PRED_HISTORY[0][24] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][24]  ( .D(\PRED_HISTORY[0][24] ), .CK(CLK), 
        .RN(n3201), .Q(\PRED_HISTORY[1][24] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][23]  ( .D(PRED[23]), .CK(CLK), .RN(n3201), .Q(
        \PRED_HISTORY[0][23] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][23]  ( .D(\PRED_HISTORY[0][23] ), .CK(CLK), 
        .RN(n3201), .Q(\PRED_HISTORY[1][23] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][22]  ( .D(PRED[22]), .CK(CLK), .RN(n3201), .Q(
        \PRED_HISTORY[0][22] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][22]  ( .D(\PRED_HISTORY[0][22] ), .CK(CLK), 
        .RN(n3201), .Q(\PRED_HISTORY[1][22] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][21]  ( .D(PRED[21]), .CK(CLK), .RN(n3201), .Q(
        \PRED_HISTORY[0][21] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][21]  ( .D(\PRED_HISTORY[0][21] ), .CK(CLK), 
        .RN(n3201), .Q(\PRED_HISTORY[1][21] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][20]  ( .D(PRED[20]), .CK(CLK), .RN(n3200), .Q(
        \PRED_HISTORY[0][20] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][20]  ( .D(\PRED_HISTORY[0][20] ), .CK(CLK), 
        .RN(n3223), .Q(\PRED_HISTORY[1][20] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][1]  ( .D(PRED[1]), .CK(CLK), .RN(n3223), .Q(
        \PRED_HISTORY[0][1] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][1]  ( .D(\PRED_HISTORY[0][1] ), .CK(CLK), .RN(
        n3223), .Q(\PRED_HISTORY[1][1] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][19]  ( .D(PRED[19]), .CK(CLK), .RN(n3223), .Q(
        \PRED_HISTORY[0][19] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][19]  ( .D(\PRED_HISTORY[0][19] ), .CK(CLK), 
        .RN(n3223), .Q(\PRED_HISTORY[1][19] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][18]  ( .D(PRED[18]), .CK(CLK), .RN(n3223), .Q(
        \PRED_HISTORY[0][18] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][18]  ( .D(\PRED_HISTORY[0][18] ), .CK(CLK), 
        .RN(n3223), .Q(\PRED_HISTORY[1][18] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][17]  ( .D(PRED[17]), .CK(CLK), .RN(n3222), .Q(
        \PRED_HISTORY[0][17] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][17]  ( .D(\PRED_HISTORY[0][17] ), .CK(CLK), 
        .RN(n3222), .Q(\PRED_HISTORY[1][17] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][16]  ( .D(PRED[16]), .CK(CLK), .RN(n3223), .Q(
        \PRED_HISTORY[0][16] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][16]  ( .D(\PRED_HISTORY[0][16] ), .CK(CLK), 
        .RN(n3223), .Q(\PRED_HISTORY[1][16] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][15]  ( .D(PRED[15]), .CK(CLK), .RN(n3223), .Q(
        \PRED_HISTORY[0][15] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][15]  ( .D(\PRED_HISTORY[0][15] ), .CK(CLK), 
        .RN(n3200), .Q(\PRED_HISTORY[1][15] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][14]  ( .D(PRED[14]), .CK(CLK), .RN(n3200), .Q(
        \PRED_HISTORY[0][14] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][14]  ( .D(\PRED_HISTORY[0][14] ), .CK(CLK), 
        .RN(n3200), .Q(\PRED_HISTORY[1][14] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][13]  ( .D(PRED[13]), .CK(CLK), .RN(n3200), .Q(
        \PRED_HISTORY[0][13] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][13]  ( .D(\PRED_HISTORY[0][13] ), .CK(CLK), 
        .RN(n3200), .Q(\PRED_HISTORY[1][13] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][12]  ( .D(PRED[12]), .CK(CLK), .RN(n3200), .Q(
        \PRED_HISTORY[0][12] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][12]  ( .D(\PRED_HISTORY[0][12] ), .CK(CLK), 
        .RN(n3200), .Q(\PRED_HISTORY[1][12] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][11]  ( .D(PRED[11]), .CK(CLK), .RN(n3200), .Q(
        \PRED_HISTORY[0][11] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][11]  ( .D(\PRED_HISTORY[0][11] ), .CK(CLK), 
        .RN(n3200), .Q(\PRED_HISTORY[1][11] ) );
  DFFR_X1 \PRED_HISTORY_reg[0][10]  ( .D(PRED[10]), .CK(CLK), .RN(n3188), .Q(
        \PRED_HISTORY[0][10] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][10]  ( .D(\PRED_HISTORY[0][10] ), .CK(CLK), 
        .RN(n3206), .Q(\PRED_HISTORY[1][10] ) );
  DFFR_X1 \PRED_HISTORY_reg[1][32]  ( .D(\PRED_HISTORY[0][32] ), .CK(CLK), 
        .RN(n3221), .Q(MISS_HIT[1]), .QN(n749) );
  DFFR_X1 \PC_HISTORY_reg[1][3]  ( .D(\PC_HISTORY[0][3] ), .CK(CLK), .RN(n3220), .QN(n750) );
  DFFR_X1 \PC_HISTORY_reg[1][2]  ( .D(\PC_HISTORY[0][2] ), .CK(CLK), .RN(n3220), .Q(n2947), .QN(n748) );
  DFFR_X1 \PC_HISTORY_reg[1][1]  ( .D(\PC_HISTORY[0][1] ), .CK(CLK), .RN(n3221), .Q(n2421), .QN(n747) );
  DFFR_X1 \PC_HISTORY_reg[1][0]  ( .D(\PC_HISTORY[0][0] ), .CK(CLK), .RN(n3220), .Q(n2946), .QN(n751) );
  DFFR_X1 \PRED_TABLE_reg[15][1]  ( .D(n1360), .CK(CLK), .RN(n3220), .Q(n2734), 
        .QN(n752) );
  DFFR_X1 \PRED_TABLE_reg[14][1]  ( .D(n1288), .CK(CLK), .RN(n3219), .Q(n2756), 
        .QN(n739) );
  DFFR_X1 \PRED_TABLE_reg[13][1]  ( .D(n1287), .CK(CLK), .RN(n3219), .Q(n2745), 
        .QN(n738) );
  DFFR_X1 \PRED_TABLE_reg[12][1]  ( .D(n1289), .CK(CLK), .RN(n3219), .Q(n2948), 
        .QN(n740) );
  DFFR_X1 \PRED_TABLE_reg[11][1]  ( .D(n1286), .CK(CLK), .RN(n3219), .Q(n2412), 
        .QN(n737) );
  DFFR_X1 \PRED_TABLE_reg[10][1]  ( .D(n1290), .CK(CLK), .RN(n3219), .Q(n2949), 
        .QN(n741) );
  DFFR_X1 \PRED_TABLE_reg[9][1]  ( .D(n1285), .CK(CLK), .RN(n3219), .Q(n2447), 
        .QN(n736) );
  DFFR_X1 \PRED_TABLE_reg[8][1]  ( .D(n1291), .CK(CLK), .RN(n3219), .QN(n742)
         );
  DFFR_X1 \PRED_TABLE_reg[7][1]  ( .D(n1284), .CK(CLK), .RN(n3220), .QN(n735)
         );
  DFFR_X1 \PRED_TABLE_reg[6][1]  ( .D(n1292), .CK(CLK), .RN(n3220), .QN(n743)
         );
  DFFR_X1 \PRED_TABLE_reg[5][1]  ( .D(n1283), .CK(CLK), .RN(n3220), .QN(n734)
         );
  DFFR_X1 \PRED_TABLE_reg[4][1]  ( .D(n1293), .CK(CLK), .RN(n3220), .Q(n2951), 
        .QN(n744) );
  DFFR_X1 \PRED_TABLE_reg[3][1]  ( .D(n1282), .CK(CLK), .RN(n3220), .QN(n733)
         );
  DFFR_X1 \PRED_TABLE_reg[2][1]  ( .D(n1294), .CK(CLK), .RN(n3220), .Q(n2767), 
        .QN(n745) );
  DFFR_X1 \PRED_TABLE_reg[1][1]  ( .D(n1281), .CK(CLK), .RN(n3220), .QN(n732)
         );
  DFFR_X1 \PRED_TABLE_reg[0][1]  ( .D(n1295), .CK(CLK), .RN(n3220), .Q(n2950), 
        .QN(n746) );
  DFFR_X1 \PC_TABLE_reg[9][5]  ( .D(n1575), .CK(CLK), .RN(n3191), .QN(n962) );
  DFFR_X1 \PC_TABLE_reg[8][5]  ( .D(n1607), .CK(CLK), .RN(n3210), .QN(n994) );
  DFFR_X1 \PC_TABLE_reg[5][2]  ( .D(n1699), .CK(CLK), .RN(n3188), .QN(n2893)
         );
  DFFR_X1 \PC_TABLE_reg[4][4]  ( .D(n1730), .CK(CLK), .RN(n3208), .Q(n418) );
  DFFR_X1 \PC_TABLE_reg[1][2]  ( .D(n1827), .CK(CLK), .RN(n3203), .Q(n390) );
  DFFR_X1 \PC_TABLE_reg[9][2]  ( .D(n1571), .CK(CLK), .RN(n3191), .QN(n958) );
  DFFR_X1 \PC_TABLE_reg[5][4]  ( .D(n1698), .CK(CLK), .RN(n3189), .QN(n2892)
         );
  DFFR_X1 \PC_TABLE_reg[10][5]  ( .D(n1543), .CK(CLK), .RN(n3215), .QN(n930)
         );
  DFFR_X1 \PC_TABLE_reg[10][3]  ( .D(n1542), .CK(CLK), .RN(n3215), .QN(n929)
         );
  DFFR_X1 \PC_TABLE_reg[3][3]  ( .D(n1766), .CK(CLK), .RN(n3233), .Q(n1961) );
  DFFR_X1 \PC_TABLE_reg[3][2]  ( .D(n1763), .CK(CLK), .RN(n3233), .Q(n1960) );
  DFFR_X1 \PC_TABLE_reg[6][4]  ( .D(n1666), .CK(CLK), .RN(n3230), .Q(n1959) );
  DFFR_X1 \PC_TABLE_reg[6][3]  ( .D(n1670), .CK(CLK), .RN(n3230), .Q(n1958) );
  DFFR_X1 \PC_TABLE_reg[12][5]  ( .D(n1479), .CK(CLK), .RN(n3199), .QN(n866)
         );
  DFFR_X1 \PC_TABLE_reg[12][4]  ( .D(n1474), .CK(CLK), .RN(n3199), .Q(n2957), 
        .QN(n861) );
  DFFR_X1 \PC_TABLE_reg[7][4]  ( .D(n1634), .CK(CLK), .RN(n3212), .QN(n2662)
         );
  DFFR_X1 \PC_TABLE_reg[7][3]  ( .D(n1638), .CK(CLK), .RN(n3212), .QN(n2789)
         );
  DFFR_X1 \PC_TABLE_reg[7][2]  ( .D(n1635), .CK(CLK), .RN(n3212), .QN(n2666)
         );
  DFFR_X1 \PC_TABLE_reg[13][5]  ( .D(n1447), .CK(CLK), .RN(n3228), .QN(n834)
         );
  DFFR_X1 \PC_TABLE_reg[13][4]  ( .D(n1442), .CK(CLK), .RN(n3228), .QN(n829)
         );
  DFFR_X1 \PC_TABLE_reg[13][2]  ( .D(n1443), .CK(CLK), .RN(n3228), .Q(n2956), 
        .QN(n830) );
  DFFR_X1 \PC_TABLE_reg[11][5]  ( .D(n1511), .CK(CLK), .RN(n3225), .QN(n898)
         );
  DFFR_X1 \PC_TABLE_reg[11][3]  ( .D(n1510), .CK(CLK), .RN(n3225), .QN(n897)
         );
  DFFR_X1 \PC_TABLE_reg[11][2]  ( .D(n1507), .CK(CLK), .RN(n3225), .QN(n894)
         );
  DFFR_X1 \PC_TABLE_reg[10][26]  ( .D(n1527), .CK(CLK), .RN(n3215), .QN(n914)
         );
  DFFR_X1 \PC_TABLE_reg[10][24]  ( .D(n1528), .CK(CLK), .RN(n3215), .QN(n915)
         );
  DFFR_X1 \PC_TABLE_reg[10][22]  ( .D(n1529), .CK(CLK), .RN(n3215), .QN(n916)
         );
  DFFR_X1 \PC_TABLE_reg[3][26]  ( .D(n1751), .CK(CLK), .RN(n3233), .Q(n1943)
         );
  DFFR_X1 \PC_TABLE_reg[3][24]  ( .D(n1752), .CK(CLK), .RN(n3233), .Q(n1942)
         );
  DFFR_X1 \PC_TABLE_reg[3][22]  ( .D(n1753), .CK(CLK), .RN(n3233), .Q(n1941)
         );
  DFFR_X1 \PC_TABLE_reg[3][20]  ( .D(n1754), .CK(CLK), .RN(n3233), .Q(n1940)
         );
  DFFR_X1 \PC_TABLE_reg[10][28]  ( .D(n1526), .CK(CLK), .RN(n3214), .QN(n913)
         );
  DFFR_X1 \PC_TABLE_reg[6][26]  ( .D(n1655), .CK(CLK), .RN(n3231), .QN(n2868)
         );
  DFFR_X1 \PC_TABLE_reg[6][24]  ( .D(n1656), .CK(CLK), .RN(n3231), .QN(n2876)
         );
  DFFR_X1 \PC_TABLE_reg[6][22]  ( .D(n1657), .CK(CLK), .RN(n3231), .QN(n2874)
         );
  DFFR_X1 \PC_TABLE_reg[6][20]  ( .D(n1658), .CK(CLK), .RN(n3230), .QN(n2875)
         );
  DFFR_X1 \PC_TABLE_reg[12][26]  ( .D(n1463), .CK(CLK), .RN(n3199), .QN(n850)
         );
  DFFR_X1 \PC_TABLE_reg[12][24]  ( .D(n1464), .CK(CLK), .RN(n3199), .QN(n851)
         );
  DFFR_X1 \PC_TABLE_reg[12][22]  ( .D(n1465), .CK(CLK), .RN(n3199), .QN(n852)
         );
  DFFR_X1 \PC_TABLE_reg[12][20]  ( .D(n1466), .CK(CLK), .RN(n3199), .QN(n853)
         );
  DFFR_X1 \PC_TABLE_reg[7][24]  ( .D(n1624), .CK(CLK), .RN(n3212), .QN(n2460)
         );
  DFFR_X1 \PC_TABLE_reg[7][22]  ( .D(n1625), .CK(CLK), .RN(n3212), .QN(n2546)
         );
  DFFR_X1 \PC_TABLE_reg[7][18]  ( .D(n1627), .CK(CLK), .RN(n3235), .QN(n2514)
         );
  DFFR_X1 \PC_TABLE_reg[7][26]  ( .D(n1623), .CK(CLK), .RN(n3212), .QN(n2557)
         );
  DFFR_X1 \PC_TABLE_reg[13][24]  ( .D(n1432), .CK(CLK), .RN(n3228), .QN(n819)
         );
  DFFR_X1 \PC_TABLE_reg[13][22]  ( .D(n1433), .CK(CLK), .RN(n3228), .QN(n820)
         );
  DFFR_X1 \PC_TABLE_reg[13][18]  ( .D(n1435), .CK(CLK), .RN(n3227), .QN(n822)
         );
  DFFR_X1 \PC_TABLE_reg[11][24]  ( .D(n1496), .CK(CLK), .RN(n3225), .QN(n883)
         );
  DFFR_X1 \PC_TABLE_reg[11][20]  ( .D(n1498), .CK(CLK), .RN(n3225), .QN(n885)
         );
  DFFR_X1 \PC_TABLE_reg[13][26]  ( .D(n1431), .CK(CLK), .RN(n3228), .QN(n818)
         );
  DFFR_X1 \PC_TABLE_reg[11][18]  ( .D(n1499), .CK(CLK), .RN(n3225), .QN(n886)
         );
  DFFR_X1 \PC_TABLE_reg[11][26]  ( .D(n1495), .CK(CLK), .RN(n3225), .QN(n882)
         );
  DFFR_X1 \PC_TABLE_reg[15][5]  ( .D(n1383), .CK(CLK), .RN(n3198), .QN(n770)
         );
  DFFR_X1 \PC_TABLE_reg[15][4]  ( .D(n1379), .CK(CLK), .RN(n3198), .Q(n2959), 
        .QN(n766) );
  DFFR_X1 \PC_TABLE_reg[15][3]  ( .D(n1382), .CK(CLK), .RN(n3198), .QN(n769)
         );
  DFFR_X1 \PC_TABLE_reg[15][2]  ( .D(n1380), .CK(CLK), .RN(n3198), .Q(n2958), 
        .QN(n767) );
  DFFR_X1 \PC_TABLE_reg[14][5]  ( .D(n1415), .CK(CLK), .RN(n3195), .QN(n802)
         );
  DFFR_X1 \PC_TABLE_reg[14][4]  ( .D(n1410), .CK(CLK), .RN(n3196), .QN(n797)
         );
  DFFR_X1 \PC_TABLE_reg[14][3]  ( .D(n1414), .CK(CLK), .RN(n3196), .Q(n2955), 
        .QN(n801) );
  DFFR_X1 \PC_TABLE_reg[2][3]  ( .D(n1798), .CK(CLK), .RN(n3217), .Q(n1918) );
  DFFR_X1 \PC_TABLE_reg[10][23]  ( .D(n1552), .CK(CLK), .RN(n3216), .QN(n939)
         );
  DFFR_X1 \PC_TABLE_reg[10][21]  ( .D(n1551), .CK(CLK), .RN(n3216), .QN(n938)
         );
  DFFR_X1 \PC_TABLE_reg[10][20]  ( .D(n1530), .CK(CLK), .RN(n3215), .QN(n917)
         );
  DFFR_X1 \PC_TABLE_reg[10][19]  ( .D(n1550), .CK(CLK), .RN(n3216), .QN(n937)
         );
  DFFR_X1 \PC_TABLE_reg[10][18]  ( .D(n1531), .CK(CLK), .RN(n3215), .QN(n918)
         );
  DFFR_X1 \PC_TABLE_reg[10][17]  ( .D(n1549), .CK(CLK), .RN(n3216), .QN(n936)
         );
  DFFR_X1 \PC_TABLE_reg[10][16]  ( .D(n1532), .CK(CLK), .RN(n3215), .QN(n919)
         );
  DFFR_X1 \PC_TABLE_reg[10][15]  ( .D(n1548), .CK(CLK), .RN(n3216), .QN(n935)
         );
  DFFR_X1 \PC_TABLE_reg[10][13]  ( .D(n1547), .CK(CLK), .RN(n3216), .QN(n934)
         );
  DFFR_X1 \PC_TABLE_reg[10][6]  ( .D(n1537), .CK(CLK), .RN(n3215), .QN(n924)
         );
  DFFR_X1 \PC_TABLE_reg[10][0]  ( .D(n1540), .CK(CLK), .RN(n3215), .QN(n927)
         );
  DFFR_X1 \PC_TABLE_reg[7][31]  ( .D(n1652), .CK(CLK), .RN(n3212), .QN(n2644)
         );
  DFFR_X1 \PC_TABLE_reg[7][28]  ( .D(n1622), .CK(CLK), .RN(n3213), .QN(n2507)
         );
  DFFR_X1 \PC_TABLE_reg[7][27]  ( .D(n1650), .CK(CLK), .RN(n3213), .QN(n2472)
         );
  DFFR_X1 \PC_TABLE_reg[7][20]  ( .D(n1626), .CK(CLK), .RN(n3213), .QN(n2458)
         );
  DFFR_X1 \PC_TABLE_reg[7][19]  ( .D(n1646), .CK(CLK), .RN(n3213), .QN(n2451)
         );
  DFFR_X1 \PC_TABLE_reg[7][17]  ( .D(n1645), .CK(CLK), .RN(n3213), .QN(n2522)
         );
  DFFR_X1 \PC_TABLE_reg[7][15]  ( .D(n1644), .CK(CLK), .RN(n3213), .QN(n2535)
         );
  DFFR_X1 \PC_TABLE_reg[7][12]  ( .D(n1630), .CK(CLK), .RN(n3213), .QN(n2623)
         );
  DFFR_X1 \PC_TABLE_reg[7][11]  ( .D(n1642), .CK(CLK), .RN(n3214), .QN(n2498)
         );
  DFFR_X1 \PC_TABLE_reg[7][8]  ( .D(n1632), .CK(CLK), .RN(n3213), .QN(n2476)
         );
  DFFR_X1 \PC_TABLE_reg[7][6]  ( .D(n1633), .CK(CLK), .RN(n3213), .QN(n2655)
         );
  DFFR_X1 \PC_TABLE_reg[7][0]  ( .D(n1636), .CK(CLK), .RN(n3213), .QN(n2513)
         );
  DFFR_X1 \PC_TABLE_reg[3][23]  ( .D(n1776), .CK(CLK), .RN(n3234), .Q(n1894)
         );
  DFFR_X1 \PC_TABLE_reg[3][21]  ( .D(n1775), .CK(CLK), .RN(n3234), .Q(n1893)
         );
  DFFR_X1 \PC_TABLE_reg[3][19]  ( .D(n1774), .CK(CLK), .RN(n3234), .Q(n1892)
         );
  DFFR_X1 \PC_TABLE_reg[3][18]  ( .D(n1755), .CK(CLK), .RN(n3234), .Q(n1891)
         );
  DFFR_X1 \PC_TABLE_reg[3][17]  ( .D(n1773), .CK(CLK), .RN(n3234), .Q(n1890)
         );
  DFFR_X1 \PC_TABLE_reg[3][16]  ( .D(n1756), .CK(CLK), .RN(n3233), .Q(n1889)
         );
  DFFR_X1 \PC_TABLE_reg[3][15]  ( .D(n1772), .CK(CLK), .RN(n3234), .Q(n1888)
         );
  DFFR_X1 \PC_TABLE_reg[3][13]  ( .D(n1771), .CK(CLK), .RN(n3234), .Q(n1887)
         );
  DFFR_X1 \PC_TABLE_reg[3][6]  ( .D(n1761), .CK(CLK), .RN(n3233), .Q(n1886) );
  DFFR_X1 \PC_TABLE_reg[3][0]  ( .D(n1764), .CK(CLK), .RN(n3233), .Q(n1885) );
  DFFR_X1 \PC_TABLE_reg[10][27]  ( .D(n1554), .CK(CLK), .RN(n3214), .QN(n941)
         );
  DFFR_X1 \PC_TABLE_reg[10][12]  ( .D(n1534), .CK(CLK), .RN(n3214), .QN(n921)
         );
  DFFR_X1 \PC_TABLE_reg[10][11]  ( .D(n1546), .CK(CLK), .RN(n3214), .QN(n933)
         );
  DFFR_X1 \PC_TABLE_reg[10][7]  ( .D(n1544), .CK(CLK), .RN(n3214), .QN(n931)
         );
  DFFR_X1 \PC_TABLE_reg[10][1]  ( .D(n1541), .CK(CLK), .RN(n3214), .QN(n928)
         );
  DFFR_X1 \PC_TABLE_reg[7][25]  ( .D(n1649), .CK(CLK), .RN(n3235), .QN(n2506)
         );
  DFFR_X1 \PC_TABLE_reg[7][21]  ( .D(n1647), .CK(CLK), .RN(n3235), .QN(n2503)
         );
  DFFR_X1 \PC_TABLE_reg[7][14]  ( .D(n1629), .CK(CLK), .RN(n3212), .QN(n2601)
         );
  DFFR_X1 \PC_TABLE_reg[7][7]  ( .D(n1640), .CK(CLK), .RN(n3218), .QN(n2457)
         );
  DFFR_X1 \PC_TABLE_reg[7][1]  ( .D(n1637), .CK(CLK), .RN(n3212), .QN(n2653)
         );
  DFFR_X1 \PC_TABLE_reg[3][28]  ( .D(n1750), .CK(CLK), .RN(n3233), .Q(n1858)
         );
  DFFR_X1 \PC_TABLE_reg[3][27]  ( .D(n1778), .CK(CLK), .RN(n3232), .Q(n1831)
         );
  DFFR_X1 \PC_TABLE_reg[3][12]  ( .D(n1758), .CK(CLK), .RN(n3233), .Q(n1830)
         );
  DFFR_X1 \PC_TABLE_reg[3][11]  ( .D(n1770), .CK(CLK), .RN(n3232), .Q(n1826)
         );
  DFFR_X1 \PC_TABLE_reg[3][7]  ( .D(n1768), .CK(CLK), .RN(n3232), .Q(n1799) );
  DFFR_X1 \PC_TABLE_reg[3][1]  ( .D(n1765), .CK(CLK), .RN(n3233), .Q(n1795) );
  DFFR_X1 \PC_TABLE_reg[10][31]  ( .D(n1556), .CK(CLK), .RN(n3215), .QN(n943)
         );
  DFFR_X1 \PC_TABLE_reg[10][30]  ( .D(n1525), .CK(CLK), .RN(n3216), .QN(n912)
         );
  DFFR_X1 \PC_TABLE_reg[10][29]  ( .D(n1555), .CK(CLK), .RN(n3216), .QN(n942)
         );
  DFFR_X1 \PC_TABLE_reg[10][25]  ( .D(n1553), .CK(CLK), .RN(n3216), .QN(n940)
         );
  DFFR_X1 \PC_TABLE_reg[10][14]  ( .D(n1533), .CK(CLK), .RN(n3216), .QN(n920)
         );
  DFFR_X1 \PC_TABLE_reg[10][10]  ( .D(n1535), .CK(CLK), .RN(n3216), .QN(n922)
         );
  DFFR_X1 \PC_TABLE_reg[10][9]  ( .D(n1545), .CK(CLK), .RN(n3216), .QN(n932)
         );
  DFFR_X1 \PC_TABLE_reg[10][8]  ( .D(n1536), .CK(CLK), .RN(n3215), .QN(n923)
         );
  DFFR_X1 \PC_TABLE_reg[7][30]  ( .D(n1621), .CK(CLK), .RN(n3214), .QN(n2568)
         );
  DFFR_X1 \PC_TABLE_reg[7][29]  ( .D(n1651), .CK(CLK), .RN(n3214), .QN(n2579)
         );
  DFFR_X1 \PC_TABLE_reg[7][23]  ( .D(n1648), .CK(CLK), .RN(n3214), .QN(n2455)
         );
  DFFR_X1 \PC_TABLE_reg[7][16]  ( .D(n1628), .CK(CLK), .RN(n3213), .QN(n2450)
         );
  DFFR_X1 \PC_TABLE_reg[7][13]  ( .D(n1643), .CK(CLK), .RN(n3214), .QN(n2612)
         );
  DFFR_X1 \PC_TABLE_reg[7][10]  ( .D(n1631), .CK(CLK), .RN(n3213), .QN(n2590)
         );
  DFFR_X1 \PC_TABLE_reg[7][9]  ( .D(n1641), .CK(CLK), .RN(n3214), .QN(n2512)
         );
  DFFR_X1 \PC_TABLE_reg[3][31]  ( .D(n1780), .CK(CLK), .RN(n3234), .Q(n1570)
         );
  DFFR_X1 \PC_TABLE_reg[3][30]  ( .D(n1749), .CK(CLK), .RN(n3235), .Q(n1539)
         );
  DFFR_X1 \PC_TABLE_reg[3][29]  ( .D(n1779), .CK(CLK), .RN(n3234), .Q(n1538)
         );
  DFFR_X1 \PC_TABLE_reg[3][25]  ( .D(n1777), .CK(CLK), .RN(n3235), .Q(n1506)
         );
  DFFR_X1 \PC_TABLE_reg[3][14]  ( .D(n1757), .CK(CLK), .RN(n3234), .Q(n1478)
         );
  DFFR_X1 \PC_TABLE_reg[3][10]  ( .D(n1759), .CK(CLK), .RN(n3234), .Q(n1475)
         );
  DFFR_X1 \PC_TABLE_reg[3][9]  ( .D(n1769), .CK(CLK), .RN(n3235), .Q(n1446) );
  DFFR_X1 \PC_TABLE_reg[3][8]  ( .D(n1760), .CK(CLK), .RN(n3234), .Q(n1411) );
  DFFR_X1 \PC_TABLE_reg[6][23]  ( .D(n1680), .CK(CLK), .RN(n3231), .QN(n2844)
         );
  DFFR_X1 \PC_TABLE_reg[6][21]  ( .D(n1679), .CK(CLK), .RN(n3232), .QN(n2822)
         );
  DFFR_X1 \PC_TABLE_reg[6][19]  ( .D(n1678), .CK(CLK), .RN(n3232), .QN(n2833)
         );
  DFFR_X1 \PC_TABLE_reg[6][18]  ( .D(n1659), .CK(CLK), .RN(n3231), .QN(n2872)
         );
  DFFR_X1 \PC_TABLE_reg[6][17]  ( .D(n1677), .CK(CLK), .RN(n3232), .QN(n2800)
         );
  DFFR_X1 \PC_TABLE_reg[6][16]  ( .D(n1660), .CK(CLK), .RN(n3231), .QN(n2867)
         );
  DFFR_X1 \PC_TABLE_reg[6][15]  ( .D(n1676), .CK(CLK), .RN(n3232), .QN(n2873)
         );
  DFFR_X1 \PC_TABLE_reg[6][13]  ( .D(n1675), .CK(CLK), .RN(n3232), .QN(n2871)
         );
  DFFR_X1 \PC_TABLE_reg[6][6]  ( .D(n1665), .CK(CLK), .RN(n3231), .QN(n2885)
         );
  DFFR_X1 \PC_TABLE_reg[6][0]  ( .D(n1668), .CK(CLK), .RN(n3231), .QN(n2866)
         );
  DFFR_X1 \PC_TABLE_reg[6][28]  ( .D(n1654), .CK(CLK), .RN(n3230), .QN(n2878)
         );
  DFFR_X1 \PC_TABLE_reg[6][27]  ( .D(n1682), .CK(CLK), .RN(n3230), .QN(n2811)
         );
  DFFR_X1 \PC_TABLE_reg[6][12]  ( .D(n1662), .CK(CLK), .RN(n3230), .QN(n2882)
         );
  DFFR_X1 \PC_TABLE_reg[6][11]  ( .D(n1674), .CK(CLK), .RN(n3230), .QN(n2883)
         );
  DFFR_X1 \PC_TABLE_reg[6][7]  ( .D(n1672), .CK(CLK), .RN(n3230), .QN(n2870)
         );
  DFFR_X1 \PC_TABLE_reg[6][1]  ( .D(n1669), .CK(CLK), .RN(n3230), .QN(n2884)
         );
  DFFR_X1 \PC_TABLE_reg[6][31]  ( .D(n1684), .CK(CLK), .RN(n3231), .QN(n2863)
         );
  DFFR_X1 \PC_TABLE_reg[6][30]  ( .D(n1653), .CK(CLK), .RN(n3232), .QN(n2877)
         );
  DFFR_X1 \PC_TABLE_reg[6][29]  ( .D(n1683), .CK(CLK), .RN(n3232), .QN(n1070)
         );
  DFFR_X1 \PC_TABLE_reg[6][25]  ( .D(n1681), .CK(CLK), .RN(n3232), .QN(n1068)
         );
  DFFR_X1 \PC_TABLE_reg[6][14]  ( .D(n1661), .CK(CLK), .RN(n3231), .QN(n2881)
         );
  DFFR_X1 \PC_TABLE_reg[6][10]  ( .D(n1663), .CK(CLK), .RN(n3231), .QN(n2869)
         );
  DFFR_X1 \PC_TABLE_reg[6][9]  ( .D(n1673), .CK(CLK), .RN(n3232), .QN(n2879)
         );
  DFFR_X1 \PC_TABLE_reg[6][8]  ( .D(n1664), .CK(CLK), .RN(n3231), .QN(n2880)
         );
  DFFR_X1 \PC_TABLE_reg[13][31]  ( .D(n1460), .CK(CLK), .RN(n3228), .QN(n2891)
         );
  DFFR_X1 \PC_TABLE_reg[13][28]  ( .D(n1430), .CK(CLK), .RN(n3229), .QN(n2889)
         );
  DFFR_X1 \PC_TABLE_reg[13][27]  ( .D(n1458), .CK(CLK), .RN(n3229), .QN(n2890)
         );
  DFFR_X1 \PC_TABLE_reg[13][20]  ( .D(n1434), .CK(CLK), .RN(n3229), .QN(n2887)
         );
  DFFR_X1 \PC_TABLE_reg[13][19]  ( .D(n1454), .CK(CLK), .RN(n3229), .QN(n2888)
         );
  DFFR_X1 \PC_TABLE_reg[13][17]  ( .D(n1453), .CK(CLK), .RN(n3229), .QN(n2886)
         );
  DFFR_X1 \PC_TABLE_reg[13][15]  ( .D(n1452), .CK(CLK), .RN(n3229), .QN(n839)
         );
  DFFR_X1 \PC_TABLE_reg[13][12]  ( .D(n1438), .CK(CLK), .RN(n3228), .QN(n825)
         );
  DFFR_X1 \PC_TABLE_reg[13][11]  ( .D(n1450), .CK(CLK), .RN(n3229), .QN(n837)
         );
  DFFR_X1 \PC_TABLE_reg[13][8]  ( .D(n1440), .CK(CLK), .RN(n3228), .QN(n827)
         );
  DFFR_X1 \PC_TABLE_reg[13][6]  ( .D(n1441), .CK(CLK), .RN(n3228), .QN(n828)
         );
  DFFR_X1 \PC_TABLE_reg[13][0]  ( .D(n1444), .CK(CLK), .RN(n3228), .QN(n831)
         );
  DFFR_X1 \PC_TABLE_reg[13][25]  ( .D(n1457), .CK(CLK), .RN(n3227), .QN(n844)
         );
  DFFR_X1 \PC_TABLE_reg[13][21]  ( .D(n1455), .CK(CLK), .RN(n3227), .QN(n842)
         );
  DFFR_X1 \PC_TABLE_reg[13][14]  ( .D(n1437), .CK(CLK), .RN(n3227), .QN(n824)
         );
  DFFR_X1 \PC_TABLE_reg[13][7]  ( .D(n1448), .CK(CLK), .RN(n3227), .QN(n835)
         );
  DFFR_X1 \PC_TABLE_reg[13][1]  ( .D(n1445), .CK(CLK), .RN(n3228), .QN(n832)
         );
  DFFR_X1 \PC_TABLE_reg[12][23]  ( .D(n1488), .CK(CLK), .RN(n3224), .QN(n875)
         );
  DFFR_X1 \PC_TABLE_reg[12][21]  ( .D(n1487), .CK(CLK), .RN(n3224), .QN(n874)
         );
  DFFR_X1 \PC_TABLE_reg[12][19]  ( .D(n1486), .CK(CLK), .RN(n3224), .QN(n873)
         );
  DFFR_X1 \PC_TABLE_reg[12][18]  ( .D(n1467), .CK(CLK), .RN(n3200), .QN(n854)
         );
  DFFR_X1 \PC_TABLE_reg[12][17]  ( .D(n1485), .CK(CLK), .RN(n3224), .QN(n872)
         );
  DFFR_X1 \PC_TABLE_reg[12][16]  ( .D(n1468), .CK(CLK), .RN(n3200), .QN(n855)
         );
  DFFR_X1 \PC_TABLE_reg[12][15]  ( .D(n1484), .CK(CLK), .RN(n3224), .QN(n871)
         );
  DFFR_X1 \PC_TABLE_reg[12][13]  ( .D(n1483), .CK(CLK), .RN(n3224), .QN(n870)
         );
  DFFR_X1 \PC_TABLE_reg[12][6]  ( .D(n1473), .CK(CLK), .RN(n3199), .QN(n860)
         );
  DFFR_X1 \PC_TABLE_reg[12][0]  ( .D(n1476), .CK(CLK), .RN(n3199), .QN(n863)
         );
  DFFR_X1 \PC_TABLE_reg[12][28]  ( .D(n1462), .CK(CLK), .RN(n3199), .QN(n849)
         );
  DFFR_X1 \PC_TABLE_reg[12][27]  ( .D(n1490), .CK(CLK), .RN(n3198), .QN(n877)
         );
  DFFR_X1 \PC_TABLE_reg[12][12]  ( .D(n1470), .CK(CLK), .RN(n3199), .QN(n857)
         );
  DFFR_X1 \PC_TABLE_reg[12][11]  ( .D(n1482), .CK(CLK), .RN(n3198), .QN(n869)
         );
  DFFR_X1 \PC_TABLE_reg[12][7]  ( .D(n1480), .CK(CLK), .RN(n3199), .QN(n867)
         );
  DFFR_X1 \PC_TABLE_reg[12][1]  ( .D(n1477), .CK(CLK), .RN(n3199), .QN(n864)
         );
  DFFR_X1 \PC_TABLE_reg[11][31]  ( .D(n1524), .CK(CLK), .RN(n3226), .QN(n911)
         );
  DFFR_X1 \PC_TABLE_reg[11][28]  ( .D(n1494), .CK(CLK), .RN(n3226), .QN(n881)
         );
  DFFR_X1 \PC_TABLE_reg[11][27]  ( .D(n1522), .CK(CLK), .RN(n3226), .QN(n909)
         );
  DFFR_X1 \PC_TABLE_reg[11][22]  ( .D(n1497), .CK(CLK), .RN(n3226), .QN(n884)
         );
  DFFR_X1 \PC_TABLE_reg[11][19]  ( .D(n1518), .CK(CLK), .RN(n3226), .QN(n905)
         );
  DFFR_X1 \PC_TABLE_reg[11][17]  ( .D(n1517), .CK(CLK), .RN(n3226), .QN(n904)
         );
  DFFR_X1 \PC_TABLE_reg[11][15]  ( .D(n1516), .CK(CLK), .RN(n3227), .QN(n903)
         );
  DFFR_X1 \PC_TABLE_reg[11][12]  ( .D(n1502), .CK(CLK), .RN(n3226), .QN(n889)
         );
  DFFR_X1 \PC_TABLE_reg[11][11]  ( .D(n1514), .CK(CLK), .RN(n3227), .QN(n901)
         );
  DFFR_X1 \PC_TABLE_reg[11][8]  ( .D(n1504), .CK(CLK), .RN(n3226), .QN(n891)
         );
  DFFR_X1 \PC_TABLE_reg[11][6]  ( .D(n1505), .CK(CLK), .RN(n3226), .QN(n892)
         );
  DFFR_X1 \PC_TABLE_reg[11][0]  ( .D(n1508), .CK(CLK), .RN(n3226), .QN(n895)
         );
  DFFR_X1 \PC_TABLE_reg[13][30]  ( .D(n1429), .CK(CLK), .RN(n3230), .QN(n816)
         );
  DFFR_X1 \PC_TABLE_reg[13][29]  ( .D(n1459), .CK(CLK), .RN(n3229), .QN(n846)
         );
  DFFR_X1 \PC_TABLE_reg[13][23]  ( .D(n1456), .CK(CLK), .RN(n3229), .QN(n843)
         );
  DFFR_X1 \PC_TABLE_reg[13][16]  ( .D(n1436), .CK(CLK), .RN(n3229), .QN(n823)
         );
  DFFR_X1 \PC_TABLE_reg[13][13]  ( .D(n1451), .CK(CLK), .RN(n3230), .QN(n838)
         );
  DFFR_X1 \PC_TABLE_reg[13][10]  ( .D(n1439), .CK(CLK), .RN(n3229), .QN(n826)
         );
  DFFR_X1 \PC_TABLE_reg[13][9]  ( .D(n1449), .CK(CLK), .RN(n3230), .QN(n836)
         );
  DFFR_X1 \PC_TABLE_reg[11][25]  ( .D(n1521), .CK(CLK), .RN(n3225), .QN(n908)
         );
  DFFR_X1 \PC_TABLE_reg[11][21]  ( .D(n1519), .CK(CLK), .RN(n3225), .QN(n906)
         );
  DFFR_X1 \PC_TABLE_reg[11][14]  ( .D(n1501), .CK(CLK), .RN(n3225), .QN(n888)
         );
  DFFR_X1 \PC_TABLE_reg[11][7]  ( .D(n1512), .CK(CLK), .RN(n3225), .QN(n899)
         );
  DFFR_X1 \PC_TABLE_reg[11][1]  ( .D(n1509), .CK(CLK), .RN(n3225), .QN(n896)
         );
  DFFR_X1 \PC_TABLE_reg[12][31]  ( .D(n1492), .CK(CLK), .RN(n3229), .QN(n879)
         );
  DFFR_X1 \PC_TABLE_reg[12][30]  ( .D(n1461), .CK(CLK), .RN(n3224), .QN(n848)
         );
  DFFR_X1 \PC_TABLE_reg[12][29]  ( .D(n1491), .CK(CLK), .RN(n3224), .QN(n878)
         );
  DFFR_X1 \PC_TABLE_reg[12][25]  ( .D(n1489), .CK(CLK), .RN(n3224), .QN(n876)
         );
  DFFR_X1 \PC_TABLE_reg[12][14]  ( .D(n1469), .CK(CLK), .RN(n3224), .QN(n856)
         );
  DFFR_X1 \PC_TABLE_reg[12][10]  ( .D(n1471), .CK(CLK), .RN(n3224), .QN(n858)
         );
  DFFR_X1 \PC_TABLE_reg[12][9]  ( .D(n1481), .CK(CLK), .RN(n3224), .QN(n868)
         );
  DFFR_X1 \PC_TABLE_reg[12][8]  ( .D(n1472), .CK(CLK), .RN(n3223), .QN(n859)
         );
  DFFR_X1 \PC_TABLE_reg[11][30]  ( .D(n1493), .CK(CLK), .RN(n3227), .QN(n880)
         );
  DFFR_X1 \PC_TABLE_reg[11][29]  ( .D(n1523), .CK(CLK), .RN(n3227), .QN(n910)
         );
  DFFR_X1 \PC_TABLE_reg[11][23]  ( .D(n1520), .CK(CLK), .RN(n3227), .QN(n907)
         );
  DFFR_X1 \PC_TABLE_reg[11][16]  ( .D(n1500), .CK(CLK), .RN(n3226), .QN(n887)
         );
  DFFR_X1 \PC_TABLE_reg[11][13]  ( .D(n1515), .CK(CLK), .RN(n3227), .QN(n902)
         );
  DFFR_X1 \PC_TABLE_reg[11][10]  ( .D(n1503), .CK(CLK), .RN(n3226), .QN(n890)
         );
  DFFR_X1 \PC_TABLE_reg[11][9]  ( .D(n1513), .CK(CLK), .RN(n3227), .QN(n900)
         );
  DFFR_X1 \PC_TABLE_reg[15][26]  ( .D(n1368), .CK(CLK), .RN(n3197), .Q(n2926), 
        .QN(n755) );
  DFFR_X1 \PC_TABLE_reg[15][24]  ( .D(n1369), .CK(CLK), .RN(n3197), .Q(n2938), 
        .QN(n756) );
  DFFR_X1 \PC_TABLE_reg[15][20]  ( .D(n1371), .CK(CLK), .RN(n3196), .Q(n2935), 
        .QN(n758) );
  DFFR_X1 \PC_TABLE_reg[15][18]  ( .D(n1372), .CK(CLK), .RN(n3196), .Q(n2922), 
        .QN(n759) );
  DFFR_X1 \PC_TABLE_reg[14][0]  ( .D(n1412), .CK(CLK), .RN(n3194), .QN(n799)
         );
  DFFR_X1 \PC_TABLE_reg[14][26]  ( .D(n1399), .CK(CLK), .RN(n3195), .QN(n786)
         );
  DFFR_X1 \PC_TABLE_reg[14][24]  ( .D(n1400), .CK(CLK), .RN(n3195), .QN(n787)
         );
  DFFR_X1 \PC_TABLE_reg[14][20]  ( .D(n1402), .CK(CLK), .RN(n3194), .QN(n789)
         );
  DFFR_X1 \PC_TABLE_reg[2][25]  ( .D(n1809), .CK(CLK), .RN(n3217), .Q(n145) );
  DFFR_X1 \PC_TABLE_reg[2][23]  ( .D(n1808), .CK(CLK), .RN(n3217), .Q(n144) );
  DFFR_X1 \PC_TABLE_reg[2][22]  ( .D(n1785), .CK(CLK), .RN(n3217), .Q(n143) );
  DFFR_X1 \PC_TABLE_reg[2][21]  ( .D(n1807), .CK(CLK), .RN(n3217), .Q(n142) );
  DFFR_X1 \PC_TABLE_reg[2][20]  ( .D(n1786), .CK(CLK), .RN(n3217), .Q(n141) );
  DFFR_X1 \PC_TABLE_reg[2][18]  ( .D(n1787), .CK(CLK), .RN(n3217), .Q(n140) );
  DFFR_X1 \PC_TABLE_reg[2][7]  ( .D(n1800), .CK(CLK), .RN(n3217), .Q(n139) );
  DFFR_X1 \PC_TABLE_reg[2][1]  ( .D(n1797), .CK(CLK), .RN(n3217), .Q(n138) );
  DFFR_X1 \PC_TABLE_reg[2][0]  ( .D(n1796), .CK(CLK), .RN(n3217), .Q(n137) );
  DFFR_X1 \PC_TABLE_reg[2][31]  ( .D(n1812), .CK(CLK), .RN(n3217), .Q(n96) );
  DFFR_X1 \PC_TABLE_reg[2][30]  ( .D(n1781), .CK(CLK), .RN(n3219), .Q(n92) );
  DFFR_X1 \PC_TABLE_reg[2][29]  ( .D(n1811), .CK(CLK), .RN(n3217), .Q(n89) );
  DFFR_X1 \PC_TABLE_reg[2][27]  ( .D(n1810), .CK(CLK), .RN(n3218), .Q(n88) );
  DFFR_X1 \PC_TABLE_reg[2][16]  ( .D(n1788), .CK(CLK), .RN(n3219), .Q(n61) );
  DFFR_X1 \PC_TABLE_reg[2][14]  ( .D(n1789), .CK(CLK), .RN(n3218), .Q(n59) );
  DFFR_X1 \PC_TABLE_reg[2][13]  ( .D(n1803), .CK(CLK), .RN(n3218), .Q(n58) );
  DFFR_X1 \PC_TABLE_reg[2][12]  ( .D(n1790), .CK(CLK), .RN(n3223), .Q(n56) );
  DFFR_X1 \PC_TABLE_reg[2][11]  ( .D(n1802), .CK(CLK), .RN(n3218), .Q(n55) );
  DFFR_X1 \PC_TABLE_reg[2][9]  ( .D(n1801), .CK(CLK), .RN(n3218), .Q(n52) );
  DFFR_X1 \PC_TABLE_reg[2][28]  ( .D(n1782), .CK(CLK), .RN(n3219), .Q(n44) );
  DFFR_X1 \PC_TABLE_reg[2][26]  ( .D(n1783), .CK(CLK), .RN(n3219), .Q(n43) );
  DFFR_X1 \PC_TABLE_reg[2][24]  ( .D(n1784), .CK(CLK), .RN(n3219), .Q(n42) );
  DFFR_X1 \PC_TABLE_reg[2][19]  ( .D(n1806), .CK(CLK), .RN(n3218), .Q(n9) );
  DFFR_X1 \PC_TABLE_reg[2][17]  ( .D(n1805), .CK(CLK), .RN(n3218), .Q(n7) );
  DFFR_X1 \PC_TABLE_reg[2][15]  ( .D(n1804), .CK(CLK), .RN(n3218), .Q(n6) );
  DFFR_X1 \PC_TABLE_reg[2][10]  ( .D(n1791), .CK(CLK), .RN(n3218), .Q(n5) );
  DFFR_X1 \PC_TABLE_reg[2][8]  ( .D(n1792), .CK(CLK), .RN(n3218), .Q(n4) );
  DFFR_X1 \PC_TABLE_reg[2][6]  ( .D(n1793), .CK(CLK), .RN(n3218), .Q(n3) );
  DFFR_X1 \PC_TABLE_reg[15][31]  ( .D(n1396), .CK(CLK), .RN(n3197), .Q(n2952), 
        .QN(n783) );
  DFFR_X1 \PC_TABLE_reg[15][30]  ( .D(n1366), .CK(CLK), .RN(n3198), .Q(n2927), 
        .QN(n753) );
  DFFR_X1 \PC_TABLE_reg[15][29]  ( .D(n1395), .CK(CLK), .RN(n3197), .Q(n2928), 
        .QN(n782) );
  DFFR_X1 \PC_TABLE_reg[15][28]  ( .D(n1367), .CK(CLK), .RN(n3198), .Q(n2940), 
        .QN(n754) );
  DFFR_X1 \PC_TABLE_reg[15][27]  ( .D(n1394), .CK(CLK), .RN(n3197), .Q(n2941), 
        .QN(n781) );
  DFFR_X1 \PC_TABLE_reg[15][25]  ( .D(n1393), .CK(CLK), .RN(n3196), .Q(n2937), 
        .QN(n780) );
  DFFR_X1 \PC_TABLE_reg[15][23]  ( .D(n1392), .CK(CLK), .RN(n3196), .Q(n2939), 
        .QN(n779) );
  DFFR_X1 \PC_TABLE_reg[15][22]  ( .D(n1370), .CK(CLK), .RN(n3196), .Q(n2925), 
        .QN(n757) );
  DFFR_X1 \PC_TABLE_reg[15][21]  ( .D(n1391), .CK(CLK), .RN(n3197), .Q(n2934), 
        .QN(n778) );
  DFFR_X1 \PC_TABLE_reg[15][19]  ( .D(n1390), .CK(CLK), .RN(n3197), .Q(n2936), 
        .QN(n777) );
  DFFR_X1 \PC_TABLE_reg[15][17]  ( .D(n1389), .CK(CLK), .RN(n3198), .Q(n2923), 
        .QN(n776) );
  DFFR_X1 \PC_TABLE_reg[15][16]  ( .D(n1373), .CK(CLK), .RN(n3196), .Q(n2933), 
        .QN(n760) );
  DFFR_X1 \PC_TABLE_reg[15][15]  ( .D(n1388), .CK(CLK), .RN(n3198), .Q(n2924), 
        .QN(n775) );
  DFFR_X1 \PC_TABLE_reg[15][14]  ( .D(n1374), .CK(CLK), .RN(n3196), .Q(n2930), 
        .QN(n761) );
  DFFR_X1 \PC_TABLE_reg[15][13]  ( .D(n1387), .CK(CLK), .RN(n3198), .Q(n2931), 
        .QN(n774) );
  DFFR_X1 \PC_TABLE_reg[15][12]  ( .D(n1375), .CK(CLK), .RN(n3196), .Q(n2932), 
        .QN(n762) );
  DFFR_X1 \PC_TABLE_reg[15][11]  ( .D(n1386), .CK(CLK), .RN(n3198), .Q(n2945), 
        .QN(n773) );
  DFFR_X1 \PC_TABLE_reg[15][10]  ( .D(n1376), .CK(CLK), .RN(n3196), .Q(n2929), 
        .QN(n763) );
  DFFR_X1 \PC_TABLE_reg[15][9]  ( .D(n1385), .CK(CLK), .RN(n3197), .Q(n2942), 
        .QN(n772) );
  DFFR_X1 \PC_TABLE_reg[15][8]  ( .D(n1377), .CK(CLK), .RN(n3196), .Q(n2943), 
        .QN(n764) );
  DFFR_X1 \PC_TABLE_reg[15][7]  ( .D(n1384), .CK(CLK), .RN(n3197), .Q(n2944), 
        .QN(n771) );
  DFFR_X1 \PC_TABLE_reg[15][6]  ( .D(n1378), .CK(CLK), .RN(n3197), .Q(n2954), 
        .QN(n765) );
  DFFR_X1 \PC_TABLE_reg[15][1]  ( .D(n1381), .CK(CLK), .RN(n3197), .Q(n2953), 
        .QN(n768) );
  DFFR_X1 \PC_TABLE_reg[15][0]  ( .D(n1877), .CK(CLK), .RN(n3197), .Q(n361) );
  DFFR_X1 \PC_TABLE_reg[14][31]  ( .D(n1428), .CK(CLK), .RN(n3194), .QN(n815)
         );
  DFFR_X1 \PC_TABLE_reg[14][30]  ( .D(n1397), .CK(CLK), .RN(n3195), .QN(n784)
         );
  DFFR_X1 \PC_TABLE_reg[14][29]  ( .D(n1427), .CK(CLK), .RN(n3195), .QN(n814)
         );
  DFFR_X1 \PC_TABLE_reg[14][28]  ( .D(n1398), .CK(CLK), .RN(n3195), .QN(n785)
         );
  DFFR_X1 \PC_TABLE_reg[14][27]  ( .D(n1426), .CK(CLK), .RN(n3195), .QN(n813)
         );
  DFFR_X1 \PC_TABLE_reg[14][25]  ( .D(n1425), .CK(CLK), .RN(n3194), .QN(n812)
         );
  DFFR_X1 \PC_TABLE_reg[14][23]  ( .D(n1424), .CK(CLK), .RN(n3195), .QN(n811)
         );
  DFFR_X1 \PC_TABLE_reg[14][22]  ( .D(n1401), .CK(CLK), .RN(n3195), .QN(n788)
         );
  DFFR_X1 \PC_TABLE_reg[14][21]  ( .D(n1423), .CK(CLK), .RN(n3194), .QN(n810)
         );
  DFFR_X1 \PC_TABLE_reg[14][19]  ( .D(n1422), .CK(CLK), .RN(n3195), .QN(n809)
         );
  DFFR_X1 \PC_TABLE_reg[14][18]  ( .D(n1403), .CK(CLK), .RN(n3194), .QN(n790)
         );
  DFFR_X1 \PC_TABLE_reg[14][17]  ( .D(n1421), .CK(CLK), .RN(n3195), .QN(n808)
         );
  DFFR_X1 \PC_TABLE_reg[14][16]  ( .D(n1404), .CK(CLK), .RN(n3193), .QN(n791)
         );
  DFFR_X1 \PC_TABLE_reg[14][15]  ( .D(n1420), .CK(CLK), .RN(n3195), .QN(n807)
         );
  DFFR_X1 \PC_TABLE_reg[14][14]  ( .D(n1405), .CK(CLK), .RN(n3221), .QN(n792)
         );
  DFFR_X1 \PC_TABLE_reg[14][13]  ( .D(n1419), .CK(CLK), .RN(n3194), .QN(n806)
         );
  DFFR_X1 \PC_TABLE_reg[14][12]  ( .D(n1406), .CK(CLK), .RN(n3193), .QN(n793)
         );
  DFFR_X1 \PC_TABLE_reg[14][11]  ( .D(n1418), .CK(CLK), .RN(n3194), .QN(n805)
         );
  DFFR_X1 \PC_TABLE_reg[14][10]  ( .D(n1407), .CK(CLK), .RN(n3193), .QN(n794)
         );
  DFFR_X1 \PC_TABLE_reg[14][9]  ( .D(n1417), .CK(CLK), .RN(n3194), .QN(n804)
         );
  DFFR_X1 \PC_TABLE_reg[14][8]  ( .D(n1408), .CK(CLK), .RN(n3193), .QN(n795)
         );
  DFFR_X1 \PC_TABLE_reg[14][7]  ( .D(n1416), .CK(CLK), .RN(n3194), .QN(n803)
         );
  DFFR_X1 \PC_TABLE_reg[14][6]  ( .D(n1409), .CK(CLK), .RN(n3193), .QN(n796)
         );
  DFFR_X1 \PC_TABLE_reg[14][1]  ( .D(n1413), .CK(CLK), .RN(n3194), .QN(n800)
         );
  DFFR_X1 \PC_TABLE_reg[9][28]  ( .D(n1558), .CK(CLK), .RN(n3191), .QN(n945)
         );
  DFFR_X1 \PC_TABLE_reg[9][26]  ( .D(n1559), .CK(CLK), .RN(n3192), .QN(n946)
         );
  DFFR_X1 \PC_TABLE_reg[9][24]  ( .D(n1560), .CK(CLK), .RN(n3192), .QN(n947)
         );
  DFFR_X1 \PC_TABLE_reg[9][22]  ( .D(n1561), .CK(CLK), .RN(n3193), .QN(n948)
         );
  DFFR_X1 \PC_TABLE_reg[9][20]  ( .D(n1562), .CK(CLK), .RN(n3193), .QN(n949)
         );
  DFFR_X1 \PC_TABLE_reg[9][18]  ( .D(n1563), .CK(CLK), .RN(n3191), .QN(n950)
         );
  DFFR_X1 \PC_TABLE_reg[5][28]  ( .D(n1686), .CK(CLK), .RN(n3188), .QN(n2905)
         );
  DFFR_X1 \PC_TABLE_reg[5][26]  ( .D(n1687), .CK(CLK), .RN(n3189), .QN(n2912)
         );
  DFFR_X1 \PC_TABLE_reg[5][24]  ( .D(n1688), .CK(CLK), .RN(n3189), .QN(n2899)
         );
  DFFR_X1 \PC_TABLE_reg[5][22]  ( .D(n1689), .CK(CLK), .RN(n3190), .QN(n2911)
         );
  DFFR_X1 \PC_TABLE_reg[5][20]  ( .D(n1690), .CK(CLK), .RN(n3190), .QN(n2898)
         );
  DFFR_X1 \PC_TABLE_reg[5][18]  ( .D(n1691), .CK(CLK), .RN(n3189), .QN(n2908)
         );
  DFFR_X1 \PC_TABLE_reg[8][28]  ( .D(n1590), .CK(CLK), .RN(n3211), .QN(n977)
         );
  DFFR_X1 \PC_TABLE_reg[8][26]  ( .D(n1591), .CK(CLK), .RN(n3210), .QN(n978)
         );
  DFFR_X1 \PC_TABLE_reg[8][24]  ( .D(n1592), .CK(CLK), .RN(n3211), .QN(n979)
         );
  DFFR_X1 \PC_TABLE_reg[8][22]  ( .D(n1593), .CK(CLK), .RN(n3211), .QN(n980)
         );
  DFFR_X1 \PC_TABLE_reg[8][20]  ( .D(n1594), .CK(CLK), .RN(n3210), .QN(n981)
         );
  DFFR_X1 \PC_TABLE_reg[8][18]  ( .D(n1595), .CK(CLK), .RN(n3211), .QN(n982)
         );
  DFFR_X1 \PC_TABLE_reg[8][16]  ( .D(n1596), .CK(CLK), .RN(n3211), .QN(n983)
         );
  DFFR_X1 \PC_TABLE_reg[4][28]  ( .D(n1718), .CK(CLK), .RN(n3209), .Q(n290) );
  DFFR_X1 \PC_TABLE_reg[4][26]  ( .D(n1719), .CK(CLK), .RN(n3208), .Q(n258) );
  DFFR_X1 \PC_TABLE_reg[4][24]  ( .D(n1720), .CK(CLK), .RN(n3209), .Q(n226) );
  DFFR_X1 \PC_TABLE_reg[4][22]  ( .D(n1721), .CK(CLK), .RN(n3208), .Q(n194) );
  DFFR_X1 \PC_TABLE_reg[4][20]  ( .D(n1722), .CK(CLK), .RN(n3208), .Q(n674) );
  DFFR_X1 \PC_TABLE_reg[4][18]  ( .D(n1723), .CK(CLK), .RN(n3209), .Q(n642) );
  DFFR_X1 \PC_TABLE_reg[4][16]  ( .D(n1724), .CK(CLK), .RN(n3209), .Q(n610) );
  DFFR_X1 \PC_TABLE_reg[1][28]  ( .D(n1814), .CK(CLK), .RN(n3204), .Q(n294) );
  DFFR_X1 \PC_TABLE_reg[1][26]  ( .D(n1815), .CK(CLK), .RN(n3203), .Q(n262) );
  DFFR_X1 \PC_TABLE_reg[1][24]  ( .D(n1816), .CK(CLK), .RN(n3204), .Q(n230) );
  DFFR_X1 \PC_TABLE_reg[1][22]  ( .D(n1817), .CK(CLK), .RN(n3203), .Q(n198) );
  DFFR_X1 \PC_TABLE_reg[1][20]  ( .D(n1818), .CK(CLK), .RN(n3203), .Q(n678) );
  DFFR_X1 \PC_TABLE_reg[1][18]  ( .D(n1819), .CK(CLK), .RN(n3204), .Q(n646) );
  DFFR_X1 \PC_TABLE_reg[1][16]  ( .D(n1820), .CK(CLK), .RN(n3204), .Q(n614) );
  DFFR_X1 \PC_TABLE_reg[8][30]  ( .D(n1589), .CK(CLK), .RN(n3188), .QN(n976)
         );
  DFFR_X1 \PC_TABLE_reg[8][29]  ( .D(n1619), .CK(CLK), .RN(n3211), .QN(n2865)
         );
  DFFR_X1 \PC_TABLE_reg[8][27]  ( .D(n1618), .CK(CLK), .RN(n3212), .QN(n2679)
         );
  DFFR_X1 \PC_TABLE_reg[8][23]  ( .D(n1616), .CK(CLK), .RN(n3211), .QN(n2712)
         );
  DFFR_X1 \PC_TABLE_reg[8][21]  ( .D(n1615), .CK(CLK), .RN(n3212), .QN(n2690)
         );
  DFFR_X1 \PC_TABLE_reg[8][19]  ( .D(n1614), .CK(CLK), .RN(n3210), .QN(n2701)
         );
  DFFR_X1 \PC_TABLE_reg[8][17]  ( .D(n1613), .CK(CLK), .RN(n3211), .QN(n2668)
         );
  DFFR_X1 \PC_TABLE_reg[8][15]  ( .D(n1612), .CK(CLK), .RN(n3212), .QN(n999)
         );
  DFFR_X1 \PC_TABLE_reg[8][11]  ( .D(n1610), .CK(CLK), .RN(n3194), .QN(n997)
         );
  DFFR_X1 \PC_TABLE_reg[4][30]  ( .D(n1717), .CK(CLK), .RN(n3209), .Q(n322) );
  DFFR_X1 \PC_TABLE_reg[4][29]  ( .D(n1747), .CK(CLK), .RN(n3209), .Q(n306) );
  DFFR_X1 \PC_TABLE_reg[4][27]  ( .D(n1746), .CK(CLK), .RN(n3209), .Q(n274) );
  DFFR_X1 \PC_TABLE_reg[4][23]  ( .D(n1744), .CK(CLK), .RN(n3209), .Q(n210) );
  DFFR_X1 \PC_TABLE_reg[4][21]  ( .D(n1743), .CK(CLK), .RN(n3209), .Q(n690) );
  DFFR_X1 \PC_TABLE_reg[4][19]  ( .D(n1742), .CK(CLK), .RN(n3208), .Q(n658) );
  DFFR_X1 \PC_TABLE_reg[4][17]  ( .D(n1741), .CK(CLK), .RN(n3208), .Q(n626) );
  DFFR_X1 \PC_TABLE_reg[4][15]  ( .D(n1740), .CK(CLK), .RN(n3209), .Q(n594) );
  DFFR_X1 \PC_TABLE_reg[4][11]  ( .D(n1738), .CK(CLK), .RN(n3209), .Q(n530) );
  DFFR_X1 \PC_TABLE_reg[1][30]  ( .D(n1813), .CK(CLK), .RN(n3205), .Q(n326) );
  DFFR_X1 \PC_TABLE_reg[1][29]  ( .D(n1843), .CK(CLK), .RN(n3204), .Q(n310) );
  DFFR_X1 \PC_TABLE_reg[1][27]  ( .D(n1842), .CK(CLK), .RN(n3204), .Q(n278) );
  DFFR_X1 \PC_TABLE_reg[1][23]  ( .D(n1840), .CK(CLK), .RN(n3204), .Q(n214) );
  DFFR_X1 \PC_TABLE_reg[1][21]  ( .D(n1839), .CK(CLK), .RN(n3204), .Q(n700) );
  DFFR_X1 \PC_TABLE_reg[1][19]  ( .D(n1838), .CK(CLK), .RN(n3203), .Q(n662) );
  DFFR_X1 \PC_TABLE_reg[1][17]  ( .D(n1837), .CK(CLK), .RN(n3203), .Q(n630) );
  DFFR_X1 \PC_TABLE_reg[1][15]  ( .D(n1836), .CK(CLK), .RN(n3204), .Q(n598) );
  DFFR_X1 \PC_TABLE_reg[1][11]  ( .D(n1834), .CK(CLK), .RN(n3205), .Q(n534) );
  DFFR_X1 \PC_TABLE_reg[9][30]  ( .D(n1557), .CK(CLK), .RN(n3192), .QN(n944)
         );
  DFFR_X1 \PC_TABLE_reg[9][29]  ( .D(n1587), .CK(CLK), .RN(n3192), .QN(n974)
         );
  DFFR_X1 \PC_TABLE_reg[9][27]  ( .D(n1586), .CK(CLK), .RN(n3191), .QN(n973)
         );
  DFFR_X1 \PC_TABLE_reg[9][25]  ( .D(n1585), .CK(CLK), .RN(n3191), .QN(n972)
         );
  DFFR_X1 \PC_TABLE_reg[9][23]  ( .D(n1584), .CK(CLK), .RN(n3193), .QN(n971)
         );
  DFFR_X1 \PC_TABLE_reg[9][21]  ( .D(n1583), .CK(CLK), .RN(n3191), .QN(n970)
         );
  DFFR_X1 \PC_TABLE_reg[9][19]  ( .D(n1582), .CK(CLK), .RN(n3193), .QN(n969)
         );
  DFFR_X1 \PC_TABLE_reg[9][17]  ( .D(n1581), .CK(CLK), .RN(n3193), .QN(n968)
         );
  DFFR_X1 \PC_TABLE_reg[9][13]  ( .D(n1579), .CK(CLK), .RN(n3192), .QN(n966)
         );
  DFFR_X1 \PC_TABLE_reg[9][11]  ( .D(n1578), .CK(CLK), .RN(n3191), .QN(n965)
         );
  DFFR_X1 \PC_TABLE_reg[5][30]  ( .D(n1685), .CK(CLK), .RN(n3190), .QN(n2913)
         );
  DFFR_X1 \PC_TABLE_reg[5][29]  ( .D(n1715), .CK(CLK), .RN(n3190), .QN(n2914)
         );
  DFFR_X1 \PC_TABLE_reg[5][27]  ( .D(n1714), .CK(CLK), .RN(n3188), .QN(n2900)
         );
  DFFR_X1 \PC_TABLE_reg[5][25]  ( .D(n1713), .CK(CLK), .RN(n3189), .QN(n2904)
         );
  DFFR_X1 \PC_TABLE_reg[5][23]  ( .D(n1712), .CK(CLK), .RN(n3190), .QN(n2896)
         );
  DFFR_X1 \PC_TABLE_reg[5][21]  ( .D(n1711), .CK(CLK), .RN(n3189), .QN(n2903)
         );
  DFFR_X1 \PC_TABLE_reg[5][19]  ( .D(n1710), .CK(CLK), .RN(n3190), .QN(n2895)
         );
  DFFR_X1 \PC_TABLE_reg[5][17]  ( .D(n1709), .CK(CLK), .RN(n3190), .QN(n2909)
         );
  DFFR_X1 \PC_TABLE_reg[5][13]  ( .D(n1707), .CK(CLK), .RN(n3190), .QN(n2917)
         );
  DFFR_X1 \PC_TABLE_reg[5][11]  ( .D(n1706), .CK(CLK), .RN(n3188), .QN(n2902)
         );
  DFFR_X1 \PC_TABLE_reg[0][30]  ( .D(n1845), .CK(CLK), .RN(n3206), .Q(n325) );
  DFFR_X1 \PC_TABLE_reg[0][29]  ( .D(n1875), .CK(CLK), .RN(n3207), .Q(n309) );
  DFFR_X1 \PC_TABLE_reg[0][28]  ( .D(n1846), .CK(CLK), .RN(n3206), .Q(n293) );
  DFFR_X1 \PC_TABLE_reg[0][27]  ( .D(n1874), .CK(CLK), .RN(n3205), .Q(n277) );
  DFFR_X1 \PC_TABLE_reg[0][26]  ( .D(n1847), .CK(CLK), .RN(n3206), .Q(n261) );
  DFFR_X1 \PC_TABLE_reg[0][25]  ( .D(n1873), .CK(CLK), .RN(n3206), .Q(n245) );
  DFFR_X1 \PC_TABLE_reg[0][24]  ( .D(n1848), .CK(CLK), .RN(n3207), .Q(n229) );
  DFFR_X1 \PC_TABLE_reg[0][23]  ( .D(n1872), .CK(CLK), .RN(n3205), .Q(n213) );
  DFFR_X1 \PC_TABLE_reg[0][22]  ( .D(n1849), .CK(CLK), .RN(n3205), .Q(n197) );
  DFFR_X1 \PC_TABLE_reg[0][21]  ( .D(n1871), .CK(CLK), .RN(n3205), .Q(n699) );
  DFFR_X1 \PC_TABLE_reg[0][20]  ( .D(n1850), .CK(CLK), .RN(n3206), .Q(n677) );
  DFFR_X1 \PC_TABLE_reg[0][19]  ( .D(n1870), .CK(CLK), .RN(n3206), .Q(n661) );
  DFFR_X1 \PC_TABLE_reg[0][18]  ( .D(n1851), .CK(CLK), .RN(n3205), .Q(n645) );
  DFFR_X1 \PC_TABLE_reg[0][16]  ( .D(n1852), .CK(CLK), .RN(n3206), .Q(n613) );
  DFFR_X1 \PC_TABLE_reg[0][15]  ( .D(n1868), .CK(CLK), .RN(n3206), .Q(n597) );
  DFFR_X1 \PC_TABLE_reg[0][14]  ( .D(n1853), .CK(CLK), .RN(n3206), .Q(n581) );
  DFFR_X1 \PC_TABLE_reg[8][0]  ( .D(n1604), .CK(CLK), .RN(n3210), .QN(n991) );
  DFFR_X1 \PC_TABLE_reg[4][0]  ( .D(n1732), .CK(CLK), .RN(n3208), .Q(n354) );
  DFFR_X1 \PC_TABLE_reg[8][31]  ( .D(n1620), .CK(CLK), .RN(n3211), .QN(n2723)
         );
  DFFR_X1 \PC_TABLE_reg[8][25]  ( .D(n1617), .CK(CLK), .RN(n3188), .QN(n2864)
         );
  DFFR_X1 \PC_TABLE_reg[8][14]  ( .D(n1597), .CK(CLK), .RN(n3188), .QN(n984)
         );
  DFFR_X1 \PC_TABLE_reg[8][13]  ( .D(n1611), .CK(CLK), .RN(n3210), .QN(n998)
         );
  DFFR_X1 \PC_TABLE_reg[8][12]  ( .D(n1598), .CK(CLK), .RN(n3188), .QN(n985)
         );
  DFFR_X1 \PC_TABLE_reg[8][10]  ( .D(n1599), .CK(CLK), .RN(n3188), .QN(n986)
         );
  DFFR_X1 \PC_TABLE_reg[8][9]  ( .D(n1609), .CK(CLK), .RN(n3188), .QN(n996) );
  DFFR_X1 \PC_TABLE_reg[8][8]  ( .D(n1600), .CK(CLK), .RN(n3211), .QN(n987) );
  DFFR_X1 \PC_TABLE_reg[8][7]  ( .D(n1608), .CK(CLK), .RN(n3210), .QN(n995) );
  DFFR_X1 \PC_TABLE_reg[8][6]  ( .D(n1601), .CK(CLK), .RN(n3211), .QN(n988) );
  DFFR_X1 \PC_TABLE_reg[4][31]  ( .D(n1748), .CK(CLK), .RN(n3208), .Q(n338) );
  DFFR_X1 \PC_TABLE_reg[4][25]  ( .D(n1745), .CK(CLK), .RN(n3210), .Q(n242) );
  DFFR_X1 \PC_TABLE_reg[4][14]  ( .D(n1725), .CK(CLK), .RN(n3210), .Q(n578) );
  DFFR_X1 \PC_TABLE_reg[4][13]  ( .D(n1739), .CK(CLK), .RN(n3208), .Q(n562) );
  DFFR_X1 \PC_TABLE_reg[4][12]  ( .D(n1726), .CK(CLK), .RN(n3210), .Q(n546) );
  DFFR_X1 \PC_TABLE_reg[4][10]  ( .D(n1727), .CK(CLK), .RN(n3210), .Q(n514) );
  DFFR_X1 \PC_TABLE_reg[4][9]  ( .D(n1737), .CK(CLK), .RN(n3210), .Q(n498) );
  DFFR_X1 \PC_TABLE_reg[4][8]  ( .D(n1728), .CK(CLK), .RN(n3208), .Q(n482) );
  DFFR_X1 \PC_TABLE_reg[4][7]  ( .D(n1736), .CK(CLK), .RN(n3208), .Q(n466) );
  DFFR_X1 \PC_TABLE_reg[4][6]  ( .D(n1729), .CK(CLK), .RN(n3208), .Q(n450) );
  DFFR_X1 \PC_TABLE_reg[8][1]  ( .D(n1605), .CK(CLK), .RN(n3211), .QN(n992) );
  DFFR_X1 \PC_TABLE_reg[4][1]  ( .D(n1733), .CK(CLK), .RN(n3209), .Q(n370) );
  DFFR_X1 \PC_TABLE_reg[1][0]  ( .D(n1828), .CK(CLK), .RN(n3203), .Q(n358) );
  DFFR_X1 \PC_TABLE_reg[1][31]  ( .D(n1844), .CK(CLK), .RN(n3203), .Q(n342) );
  DFFR_X1 \PC_TABLE_reg[1][25]  ( .D(n1841), .CK(CLK), .RN(n3205), .Q(n246) );
  DFFR_X1 \PC_TABLE_reg[1][14]  ( .D(n1821), .CK(CLK), .RN(n3205), .Q(n582) );
  DFFR_X1 \PC_TABLE_reg[1][13]  ( .D(n1835), .CK(CLK), .RN(n3203), .Q(n566) );
  DFFR_X1 \PC_TABLE_reg[1][12]  ( .D(n1822), .CK(CLK), .RN(n3205), .Q(n550) );
  DFFR_X1 \PC_TABLE_reg[1][10]  ( .D(n1823), .CK(CLK), .RN(n3205), .Q(n518) );
  DFFR_X1 \PC_TABLE_reg[1][9]  ( .D(n1833), .CK(CLK), .RN(n3205), .Q(n502) );
  DFFR_X1 \PC_TABLE_reg[1][8]  ( .D(n1824), .CK(CLK), .RN(n3204), .Q(n486) );
  DFFR_X1 \PC_TABLE_reg[1][7]  ( .D(n1832), .CK(CLK), .RN(n3203), .Q(n470) );
  DFFR_X1 \PC_TABLE_reg[1][6]  ( .D(n1825), .CK(CLK), .RN(n3204), .Q(n454) );
  DFFR_X1 \PC_TABLE_reg[1][1]  ( .D(n1829), .CK(CLK), .RN(n3204), .Q(n374) );
  DFFR_X1 \PC_TABLE_reg[9][0]  ( .D(n1572), .CK(CLK), .RN(n3193), .QN(n959) );
  DFFR_X1 \PC_TABLE_reg[5][0]  ( .D(n1700), .CK(CLK), .RN(n3190), .QN(n2907)
         );
  DFFR_X1 \PC_TABLE_reg[9][31]  ( .D(n1588), .CK(CLK), .RN(n3192), .QN(n975)
         );
  DFFR_X1 \PC_TABLE_reg[9][16]  ( .D(n1564), .CK(CLK), .RN(n3193), .QN(n951)
         );
  DFFR_X1 \PC_TABLE_reg[9][15]  ( .D(n1580), .CK(CLK), .RN(n3192), .QN(n967)
         );
  DFFR_X1 \PC_TABLE_reg[9][14]  ( .D(n1565), .CK(CLK), .RN(n3192), .QN(n952)
         );
  DFFR_X1 \PC_TABLE_reg[9][12]  ( .D(n1566), .CK(CLK), .RN(n3191), .QN(n953)
         );
  DFFR_X1 \PC_TABLE_reg[9][10]  ( .D(n1567), .CK(CLK), .RN(n3192), .QN(n954)
         );
  DFFR_X1 \PC_TABLE_reg[9][9]  ( .D(n1577), .CK(CLK), .RN(n3192), .QN(n964) );
  DFFR_X1 \PC_TABLE_reg[9][8]  ( .D(n1568), .CK(CLK), .RN(n3192), .QN(n955) );
  DFFR_X1 \PC_TABLE_reg[9][7]  ( .D(n1576), .CK(CLK), .RN(n3191), .QN(n963) );
  DFFR_X1 \PC_TABLE_reg[9][6]  ( .D(n1569), .CK(CLK), .RN(n3191), .QN(n956) );
  DFFR_X1 \PC_TABLE_reg[5][31]  ( .D(n1716), .CK(CLK), .RN(n3189), .QN(n2919)
         );
  DFFR_X1 \PC_TABLE_reg[5][16]  ( .D(n1692), .CK(CLK), .RN(n3191), .QN(n2894)
         );
  DFFR_X1 \PC_TABLE_reg[5][15]  ( .D(n1708), .CK(CLK), .RN(n3190), .QN(n2910)
         );
  DFFR_X1 \PC_TABLE_reg[5][14]  ( .D(n1693), .CK(CLK), .RN(n3189), .QN(n2916)
         );
  DFFR_X1 \PC_TABLE_reg[5][12]  ( .D(n1694), .CK(CLK), .RN(n3189), .QN(n2918)
         );
  DFFR_X1 \PC_TABLE_reg[5][10]  ( .D(n1695), .CK(CLK), .RN(n3190), .QN(n2915)
         );
  DFFR_X1 \PC_TABLE_reg[5][9]  ( .D(n1705), .CK(CLK), .RN(n3190), .QN(n2906)
         );
  DFFR_X1 \PC_TABLE_reg[5][8]  ( .D(n1696), .CK(CLK), .RN(n3189), .QN(n2901)
         );
  DFFR_X1 \PC_TABLE_reg[5][7]  ( .D(n1704), .CK(CLK), .RN(n3188), .QN(n2897)
         );
  DFFR_X1 \PC_TABLE_reg[5][6]  ( .D(n1697), .CK(CLK), .RN(n3189), .QN(n2921)
         );
  DFFR_X1 \PC_TABLE_reg[9][1]  ( .D(n1573), .CK(CLK), .RN(n3192), .QN(n960) );
  DFFR_X1 \PC_TABLE_reg[5][1]  ( .D(n1701), .CK(CLK), .RN(n3189), .QN(n2920)
         );
  DFFR_X1 \PC_TABLE_reg[0][0]  ( .D(n1860), .CK(CLK), .RN(n3207), .Q(n357) );
  DFFR_X1 \PC_TABLE_reg[0][31]  ( .D(n1876), .CK(CLK), .RN(n3207), .Q(n341) );
  DFFR_X1 \PC_TABLE_reg[0][17]  ( .D(n1869), .CK(CLK), .RN(n3207), .Q(n629) );
  DFFR_X1 \PC_TABLE_reg[0][13]  ( .D(n1867), .CK(CLK), .RN(n3206), .Q(n565) );
  DFFR_X1 \PC_TABLE_reg[0][12]  ( .D(n1854), .CK(CLK), .RN(n3207), .Q(n549) );
  DFFR_X1 \PC_TABLE_reg[0][11]  ( .D(n1866), .CK(CLK), .RN(n3206), .Q(n533) );
  DFFR_X1 \PC_TABLE_reg[0][10]  ( .D(n1855), .CK(CLK), .RN(n3207), .Q(n517) );
  DFFR_X1 \PC_TABLE_reg[0][9]  ( .D(n1865), .CK(CLK), .RN(n3207), .Q(n501) );
  DFFR_X1 \PC_TABLE_reg[0][8]  ( .D(n1856), .CK(CLK), .RN(n3207), .Q(n485) );
  DFFR_X1 \PC_TABLE_reg[0][7]  ( .D(n1864), .CK(CLK), .RN(n3207), .Q(n469) );
  DFFR_X1 \PC_TABLE_reg[0][6]  ( .D(n1857), .CK(CLK), .RN(n3207), .Q(n453) );
  DFFR_X1 \PC_TABLE_reg[0][1]  ( .D(n1861), .CK(CLK), .RN(n3207), .Q(n373) );
  INV_X2 U64 ( .A(n2052), .ZN(n2053) );
  INV_X2 U123 ( .A(n3165), .ZN(n2084) );
  INV_X2 U182 ( .A(n2117), .ZN(n2116) );
  INV_X2 U242 ( .A(n3158), .ZN(n2148) );
  INV_X2 U301 ( .A(n2178), .ZN(n2179) );
  INV_X2 U365 ( .A(n3147), .ZN(n2270) );
  INV_X2 U429 ( .A(n3137), .ZN(n2335) );
  NAND3_X1 U1396 ( .A1(INST_28), .A2(n2516), .A3(n2517), .ZN(n2496) );
  BP_NB32_BP_LEN4_DW01_cmp6_0 eq_100 ( .A({\PRED_HISTORY[1][31] , 
        \PRED_HISTORY[1][30] , \PRED_HISTORY[1][29] , \PRED_HISTORY[1][28] , 
        \PRED_HISTORY[1][27] , \PRED_HISTORY[1][26] , \PRED_HISTORY[1][25] , 
        \PRED_HISTORY[1][24] , \PRED_HISTORY[1][23] , \PRED_HISTORY[1][22] , 
        \PRED_HISTORY[1][21] , \PRED_HISTORY[1][20] , \PRED_HISTORY[1][19] , 
        \PRED_HISTORY[1][18] , \PRED_HISTORY[1][17] , \PRED_HISTORY[1][16] , 
        \PRED_HISTORY[1][15] , \PRED_HISTORY[1][14] , \PRED_HISTORY[1][13] , 
        \PRED_HISTORY[1][12] , \PRED_HISTORY[1][11] , \PRED_HISTORY[1][10] , 
        \PRED_HISTORY[1][9] , \PRED_HISTORY[1][8] , \PRED_HISTORY[1][7] , 
        \PRED_HISTORY[1][6] , \PRED_HISTORY[1][5] , \PRED_HISTORY[1][4] , 
        \PRED_HISTORY[1][3] , \PRED_HISTORY[1][2] , \PRED_HISTORY[1][1] , 
        \PRED_HISTORY[1][0] }), .B(EX_PC), .TC(1'b0), .EQ(N815) );
  BP_NB32_BP_LEN4_DW01_cmp6_1 eq_59 ( .A({N90, N91, N92, N93, N94, N95, N96, 
        N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, 
        N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, 
        N121}), .B(CURR_PC), .TC(1'b0), .EQ(N122) );
  BP_NB32_BP_LEN4_DW01_add_1 add_49_2 ( .A(NEXT_PC), .B({n3182, n3182, n3182, 
        n3182, n3182, n3182, n3182, n3182, n3182, n3182, n3182, n3182, n3182, 
        n3182, n3182, n3182, n3182, INST[14:0]}), .CI(1'b0), .SUM(PRED_TK) );
  DFFS_X1 \PRED_TABLE_reg[15][0]  ( .D(n1265), .CK(CLK), .SN(n2246), .Q(n2438), 
        .QN(n716) );
  DFFS_X1 \PRED_TABLE_reg[14][0]  ( .D(n1273), .CK(CLK), .SN(n2246), .Q(n2441), 
        .QN(n724) );
  DFFS_X1 \PRED_TABLE_reg[13][0]  ( .D(n1272), .CK(CLK), .SN(n2246), .Q(n2430), 
        .QN(n723) );
  DFFS_X1 \PRED_TABLE_reg[12][0]  ( .D(n1274), .CK(CLK), .SN(n2246), .Q(n2433), 
        .QN(n725) );
  DFFS_X1 \PRED_TABLE_reg[10][0]  ( .D(n1275), .CK(CLK), .SN(n2246), .Q(n2440), 
        .QN(n726) );
  DFFS_X1 \PRED_TABLE_reg[9][0]  ( .D(n1270), .CK(CLK), .SN(n2246), .Q(n2429), 
        .QN(n721) );
  DFFS_X1 \PRED_TABLE_reg[8][0]  ( .D(n1276), .CK(CLK), .SN(n2246), .Q(n2432), 
        .QN(n727) );
  DFFS_X1 \PRED_TABLE_reg[7][0]  ( .D(n1269), .CK(CLK), .SN(n2246), .QN(n720)
         );
  DFFS_X1 \PRED_TABLE_reg[6][0]  ( .D(n1277), .CK(CLK), .SN(n2246), .QN(n728)
         );
  DFFS_X1 \PRED_TABLE_reg[5][0]  ( .D(n1268), .CK(CLK), .SN(n2246), .QN(n719)
         );
  DFFS_X1 \PRED_TABLE_reg[4][0]  ( .D(n1278), .CK(CLK), .SN(n2246), .QN(n729)
         );
  DFFS_X1 \PRED_TABLE_reg[3][0]  ( .D(n1267), .CK(CLK), .SN(n2246), .QN(n718)
         );
  DFFS_X1 \PRED_TABLE_reg[2][0]  ( .D(n1279), .CK(CLK), .SN(n2246), .QN(n730)
         );
  DFFS_X1 \PRED_TABLE_reg[1][0]  ( .D(n1266), .CK(CLK), .SN(n2246), .QN(n717)
         );
  DFFS_X1 \PRED_TABLE_reg[0][0]  ( .D(n1280), .CK(CLK), .SN(n2246), .QN(n731)
         );
  DFFS_X1 \PRED_TABLE_reg[11][0]  ( .D(n1271), .CK(CLK), .SN(n2246), .Q(n2437), 
        .QN(n722) );
  NOR2_X1 U6 ( .A1(n2855), .A2(CURR_PC[5]), .ZN(n2846) );
  NOR2_X1 U7 ( .A1(n2861), .A2(CURR_PC[2]), .ZN(n2854) );
  NOR2_X1 U8 ( .A1(n2860), .A2(CURR_PC[4]), .ZN(n2853) );
  NOR2_X1 U9 ( .A1(CURR_PC[2]), .A2(CURR_PC[3]), .ZN(n2850) );
  NAND3_X1 U10 ( .A1(n2968), .A2(n2969), .A3(n2970), .ZN(PRED[27]) );
  AND3_X1 U11 ( .A1(n2362), .A2(n2497), .A3(N122), .ZN(n3092) );
  NAND2_X1 U12 ( .A1(N815), .A2(MISS_HIT[1]), .ZN(n2407) );
  NOR2_X1 U13 ( .A1(n750), .A2(n748), .ZN(n2420) );
  NOR2_X1 U14 ( .A1(n2947), .A2(n750), .ZN(n2419) );
  NAND2_X1 U15 ( .A1(PRED_TK[27]), .A2(n3092), .ZN(n2968) );
  NAND2_X1 U16 ( .A1(NEXT_PC[27]), .A2(n3095), .ZN(n2969) );
  NAND2_X1 U17 ( .A1(NEW_PC[27]), .A2(n3105), .ZN(n2970) );
  BUF_X1 U18 ( .A(n2350), .Z(n2981) );
  BUF_X1 U19 ( .A(n2350), .Z(n2982) );
  BUF_X1 U20 ( .A(n2345), .Z(n2987) );
  BUF_X1 U21 ( .A(n2345), .Z(n2988) );
  BUF_X1 U22 ( .A(n2350), .Z(n2983) );
  BUF_X1 U23 ( .A(n2345), .Z(n2989) );
  BUF_X1 U24 ( .A(n2369), .Z(n2972) );
  BUF_X1 U25 ( .A(n2356), .Z(n2975) );
  BUF_X1 U26 ( .A(n2353), .Z(n2978) );
  BUF_X1 U27 ( .A(n2369), .Z(n2973) );
  BUF_X1 U28 ( .A(n2353), .Z(n2979) );
  BUF_X1 U29 ( .A(n2356), .Z(n2976) );
  INV_X1 U30 ( .A(n3181), .ZN(n3172) );
  INV_X1 U31 ( .A(n3181), .ZN(n3173) );
  BUF_X1 U32 ( .A(n2369), .Z(n2974) );
  BUF_X1 U33 ( .A(n2356), .Z(n2977) );
  BUF_X1 U34 ( .A(n2353), .Z(n2980) );
  INV_X1 U35 ( .A(n3134), .ZN(n2345) );
  INV_X1 U36 ( .A(n3124), .ZN(n2350) );
  BUF_X1 U37 ( .A(n2299), .Z(n2990) );
  BUF_X1 U38 ( .A(n2347), .Z(n2984) );
  BUF_X1 U39 ( .A(n2299), .Z(n2991) );
  BUF_X1 U40 ( .A(n2347), .Z(n2985) );
  BUF_X1 U41 ( .A(n2211), .Z(n2993) );
  BUF_X1 U42 ( .A(n2211), .Z(n2994) );
  BUF_X1 U43 ( .A(n2299), .Z(n2992) );
  BUF_X1 U44 ( .A(n2344), .Z(n3131) );
  BUF_X1 U45 ( .A(n2344), .Z(n3133) );
  BUF_X1 U46 ( .A(n2344), .Z(n3132) );
  BUF_X1 U47 ( .A(n2344), .Z(n3134) );
  BUF_X1 U48 ( .A(n2347), .Z(n2986) );
  BUF_X1 U49 ( .A(n2351), .Z(n3121) );
  BUF_X1 U50 ( .A(n2351), .Z(n3122) );
  BUF_X1 U51 ( .A(n2351), .Z(n3123) );
  BUF_X1 U52 ( .A(n2351), .Z(n3124) );
  BUF_X1 U53 ( .A(n2211), .Z(n2995) );
  BUF_X1 U54 ( .A(n2344), .Z(n3135) );
  BUF_X1 U55 ( .A(n2351), .Z(n3125) );
  BUF_X1 U56 ( .A(n3171), .Z(n3181) );
  BUF_X1 U57 ( .A(n3169), .Z(n3176) );
  BUF_X1 U58 ( .A(n3170), .Z(n3178) );
  BUF_X1 U59 ( .A(n3170), .Z(n3177) );
  BUF_X1 U60 ( .A(n3169), .Z(n3175) );
  BUF_X1 U61 ( .A(n3169), .Z(n3174) );
  BUF_X1 U62 ( .A(n3170), .Z(n3179) );
  BUF_X1 U63 ( .A(n3171), .Z(n3180) );
  INV_X1 U65 ( .A(n3109), .ZN(n2369) );
  INV_X1 U66 ( .A(n3119), .ZN(n2353) );
  INV_X1 U67 ( .A(n3114), .ZN(n2356) );
  NOR2_X1 U68 ( .A1(n3010), .A2(n2114), .ZN(n2344) );
  NOR2_X1 U69 ( .A1(n3003), .A2(n2114), .ZN(n2351) );
  BUF_X1 U70 ( .A(n2271), .Z(n3146) );
  BUF_X1 U71 ( .A(n2271), .Z(n3147) );
  BUF_X1 U72 ( .A(n2271), .Z(n3148) );
  BUF_X1 U73 ( .A(n2271), .Z(n3149) );
  BUF_X1 U74 ( .A(n2370), .Z(n3106) );
  BUF_X1 U75 ( .A(n2370), .Z(n3108) );
  BUF_X1 U76 ( .A(n2370), .Z(n3107) );
  BUF_X1 U77 ( .A(n2354), .Z(n3117) );
  BUF_X1 U78 ( .A(n2354), .Z(n3116) );
  BUF_X1 U79 ( .A(n2354), .Z(n3118) );
  BUF_X1 U80 ( .A(n2370), .Z(n3109) );
  BUF_X1 U81 ( .A(n2354), .Z(n3119) );
  BUF_X1 U82 ( .A(n2357), .Z(n3113) );
  BUF_X1 U83 ( .A(n2357), .Z(n3112) );
  BUF_X1 U84 ( .A(n2357), .Z(n3111) );
  BUF_X1 U85 ( .A(n2357), .Z(n3114) );
  BUF_X1 U86 ( .A(n2370), .Z(n3110) );
  BUF_X1 U87 ( .A(n2354), .Z(n3120) );
  BUF_X1 U88 ( .A(n2357), .Z(n3115) );
  INV_X1 U89 ( .A(n3129), .ZN(n2347) );
  INV_X1 U90 ( .A(n3141), .ZN(n2299) );
  INV_X1 U91 ( .A(n3150), .ZN(n2211) );
  BUF_X1 U92 ( .A(n2049), .Z(n3169) );
  BUF_X1 U93 ( .A(n2049), .Z(n3170) );
  BUF_X1 U94 ( .A(n2049), .Z(n3171) );
  INV_X1 U95 ( .A(n2082), .ZN(n2114) );
  NOR2_X1 U96 ( .A1(n3023), .A2(n2114), .ZN(n2370) );
  NOR2_X1 U97 ( .A1(n3029), .A2(n2114), .ZN(n2357) );
  NOR2_X1 U98 ( .A1(n3046), .A2(n2114), .ZN(n2354) );
  BUF_X1 U99 ( .A(n2147), .Z(n3159) );
  BUF_X1 U100 ( .A(n2147), .Z(n3158) );
  BUF_X1 U101 ( .A(n2085), .Z(n3164) );
  NOR2_X1 U102 ( .A1(n3079), .A2(n2114), .ZN(n2271) );
  BUF_X1 U103 ( .A(n2147), .Z(n3160) );
  BUF_X1 U104 ( .A(n2085), .Z(n3166) );
  BUF_X1 U105 ( .A(n2085), .Z(n3165) );
  NOR2_X1 U106 ( .A1(n2372), .A2(n2114), .ZN(n2049) );
  BUF_X1 U107 ( .A(n2147), .Z(n3157) );
  BUF_X1 U108 ( .A(n2085), .Z(n3163) );
  BUF_X1 U109 ( .A(n2333), .Z(n3136) );
  BUF_X1 U110 ( .A(n2348), .Z(n3126) );
  BUF_X1 U111 ( .A(n2348), .Z(n3127) );
  BUF_X1 U112 ( .A(n2348), .Z(n3128) );
  BUF_X1 U113 ( .A(n2333), .Z(n3137) );
  BUF_X1 U114 ( .A(n2348), .Z(n3129) );
  BUF_X1 U115 ( .A(n2333), .Z(n3138) );
  BUF_X1 U116 ( .A(n2333), .Z(n3139) );
  BUF_X1 U117 ( .A(n2300), .Z(n3141) );
  BUF_X1 U118 ( .A(n2300), .Z(n3143) );
  BUF_X1 U119 ( .A(n2300), .Z(n3144) );
  BUF_X1 U120 ( .A(n2300), .Z(n3142) );
  BUF_X1 U121 ( .A(n2208), .Z(n3150) );
  BUF_X1 U122 ( .A(n2208), .Z(n3151) );
  BUF_X1 U124 ( .A(n2208), .Z(n3153) );
  BUF_X1 U125 ( .A(n2208), .Z(n3152) );
  NAND2_X1 U126 ( .A1(n3059), .A2(n2082), .ZN(n2178) );
  NAND2_X1 U127 ( .A1(n3077), .A2(n2082), .ZN(n2117) );
  BUF_X1 U128 ( .A(n2333), .Z(n3140) );
  BUF_X1 U129 ( .A(n2348), .Z(n3130) );
  BUF_X1 U130 ( .A(n2300), .Z(n3145) );
  BUF_X1 U131 ( .A(n2208), .Z(n3154) );
  INV_X2 U132 ( .A(n2372), .ZN(n2504) );
  INV_X1 U133 ( .A(n3082), .ZN(n2659) );
  INV_X1 U134 ( .A(n3047), .ZN(n2509) );
  INV_X1 U135 ( .A(n3030), .ZN(n2510) );
  INV_X1 U136 ( .A(n3024), .ZN(n2661) );
  BUF_X1 U137 ( .A(n3187), .Z(n3244) );
  BUF_X1 U138 ( .A(n3183), .Z(n3237) );
  BUF_X1 U139 ( .A(n3185), .Z(n3240) );
  BUF_X1 U140 ( .A(n3185), .Z(n3241) );
  BUF_X1 U141 ( .A(n3183), .Z(n3236) );
  BUF_X1 U142 ( .A(n3184), .Z(n3238) );
  BUF_X1 U143 ( .A(n3186), .Z(n3243) );
  BUF_X1 U144 ( .A(n3184), .Z(n3239) );
  BUF_X1 U145 ( .A(n3186), .Z(n3242) );
  BUF_X1 U146 ( .A(n3187), .Z(n3245) );
  BUF_X1 U147 ( .A(n2463), .Z(n3094) );
  AND3_X1 U148 ( .A1(n2362), .A2(n2497), .A3(N122), .ZN(n3091) );
  NOR2_X1 U149 ( .A1(n2496), .A2(N122), .ZN(n2082) );
  NOR2_X1 U150 ( .A1(n3018), .A2(n2114), .ZN(n2348) );
  NOR2_X1 U151 ( .A1(n3090), .A2(n2114), .ZN(n2300) );
  NOR2_X1 U152 ( .A1(n3087), .A2(n2114), .ZN(n2208) );
  NOR2_X1 U153 ( .A1(n3083), .A2(n2114), .ZN(n2333) );
  NOR2_X1 U154 ( .A1(n2113), .A2(n2114), .ZN(n2085) );
  INV_X1 U155 ( .A(n2496), .ZN(n2362) );
  NOR2_X1 U156 ( .A1(n2176), .A2(n2114), .ZN(n2147) );
  BUF_X1 U157 ( .A(n2463), .Z(n3093) );
  AND3_X1 U158 ( .A1(n2362), .A2(n2497), .A3(N122), .ZN(n2462) );
  BUF_X1 U159 ( .A(n2463), .Z(n3095) );
  NAND2_X1 U160 ( .A1(n3085), .A2(n2082), .ZN(n2052) );
  NOR2_X1 U161 ( .A1(n2362), .A2(n2408), .ZN(n2464) );
  NOR2_X1 U162 ( .A1(n2362), .A2(n2408), .ZN(n3097) );
  NOR2_X1 U163 ( .A1(n2362), .A2(n2408), .ZN(n3096) );
  INV_X2 U164 ( .A(n2113), .ZN(n2526) );
  INV_X2 U165 ( .A(n2176), .ZN(n2525) );
  NAND2_X1 U166 ( .A1(n2847), .A2(n2849), .ZN(n2372) );
  BUF_X1 U167 ( .A(n2298), .Z(n3079) );
  BUF_X1 U168 ( .A(n2298), .Z(n3080) );
  BUF_X1 U169 ( .A(n2298), .Z(n3081) );
  INV_X1 U170 ( .A(n2352), .ZN(n2999) );
  INV_X1 U171 ( .A(n2352), .ZN(n3001) );
  INV_X1 U172 ( .A(n2346), .ZN(n3009) );
  INV_X1 U173 ( .A(n2352), .ZN(n3000) );
  INV_X1 U174 ( .A(n2346), .ZN(n3008) );
  BUF_X1 U175 ( .A(n2298), .Z(n3082) );
  BUF_X1 U176 ( .A(n3026), .Z(n3027) );
  BUF_X1 U177 ( .A(n3026), .Z(n3028) );
  BUF_X1 U178 ( .A(n3019), .Z(n3020) );
  BUF_X1 U179 ( .A(n3019), .Z(n3022) );
  BUF_X1 U180 ( .A(n3019), .Z(n3021) );
  BUF_X1 U181 ( .A(n3049), .Z(n3051) );
  BUF_X1 U183 ( .A(n3050), .Z(n3055) );
  BUF_X1 U184 ( .A(n3050), .Z(n3056) );
  BUF_X1 U185 ( .A(n3050), .Z(n3057) );
  BUF_X1 U186 ( .A(n3049), .Z(n3052) );
  BUF_X1 U187 ( .A(n3049), .Z(n3054) );
  BUF_X1 U188 ( .A(n3049), .Z(n3053) );
  BUF_X1 U189 ( .A(n3026), .Z(n3029) );
  BUF_X1 U190 ( .A(n2368), .Z(n3030) );
  BUF_X1 U191 ( .A(n2371), .Z(n3023) );
  BUF_X1 U192 ( .A(n2371), .Z(n3024) );
  BUF_X1 U193 ( .A(n2371), .Z(n3025) );
  BUF_X1 U194 ( .A(n2368), .Z(n3032) );
  BUF_X1 U195 ( .A(n2368), .Z(n3031) );
  BUF_X1 U196 ( .A(n3050), .Z(n3058) );
  BUF_X1 U197 ( .A(n2207), .Z(n3060) );
  BUF_X1 U198 ( .A(n2207), .Z(n3061) );
  BUF_X1 U199 ( .A(n2207), .Z(n3062) );
  BUF_X1 U200 ( .A(n2207), .Z(n3059) );
  INV_X1 U201 ( .A(n2375), .ZN(n2373) );
  INV_X1 U202 ( .A(n2405), .ZN(n2404) );
  INV_X1 U203 ( .A(n2401), .ZN(n2400) );
  INV_X1 U204 ( .A(n2397), .ZN(n2396) );
  INV_X1 U205 ( .A(n2393), .ZN(n2392) );
  INV_X1 U206 ( .A(n2391), .ZN(n2390) );
  INV_X1 U207 ( .A(n2389), .ZN(n2388) );
  INV_X1 U208 ( .A(n2387), .ZN(n2386) );
  INV_X1 U209 ( .A(n2385), .ZN(n2384) );
  INV_X1 U210 ( .A(n2383), .ZN(n2382) );
  INV_X1 U211 ( .A(n2381), .ZN(n2380) );
  INV_X1 U212 ( .A(n2379), .ZN(n2378) );
  INV_X1 U213 ( .A(n2377), .ZN(n2376) );
  INV_X1 U214 ( .A(n2395), .ZN(n2394) );
  INV_X1 U215 ( .A(n2403), .ZN(n2402) );
  INV_X1 U216 ( .A(n2399), .ZN(n2398) );
  INV_X1 U217 ( .A(n2482), .ZN(PRED[21]) );
  AOI222_X1 U218 ( .A1(PRED_TK[21]), .A2(n3092), .B1(NEXT_PC[21]), .B2(n3094), 
        .C1(NEW_PC[21]), .C2(n3104), .ZN(n2482) );
  INV_X1 U219 ( .A(n2461), .ZN(PRED[9]) );
  AOI222_X1 U220 ( .A1(PRED_TK[9]), .A2(n3092), .B1(NEXT_PC[9]), .B2(n3094), 
        .C1(NEW_PC[9]), .C2(n3102), .ZN(n2461) );
  INV_X1 U221 ( .A(n2407), .ZN(n2408) );
  OAI22_X1 U222 ( .A1(n3139), .A2(n2864), .B1(n2217), .B2(n2335), .ZN(n1617)
         );
  OAI22_X1 U223 ( .A1(n3139), .A2(n2723), .B1(n2210), .B2(n2335), .ZN(n1620)
         );
  OAI22_X1 U224 ( .A1(n3139), .A2(n2668), .B1(n2225), .B2(n2335), .ZN(n1613)
         );
  OAI22_X1 U225 ( .A1(n3140), .A2(n2701), .B1(n2223), .B2(n2335), .ZN(n1614)
         );
  OAI22_X1 U226 ( .A1(n3136), .A2(n2690), .B1(n2221), .B2(n2335), .ZN(n1615)
         );
  OAI22_X1 U227 ( .A1(n3138), .A2(n2712), .B1(n2219), .B2(n2335), .ZN(n1616)
         );
  OAI22_X1 U228 ( .A1(n3137), .A2(n2679), .B1(n2215), .B2(n2335), .ZN(n1618)
         );
  OAI22_X1 U229 ( .A1(n3138), .A2(n2865), .B1(n2213), .B2(n2335), .ZN(n1619)
         );
  INV_X1 U230 ( .A(INST_27), .ZN(n2516) );
  NOR3_X1 U231 ( .A1(INST_29), .A2(INST_31), .A3(INST_30), .ZN(n2517) );
  OAI22_X1 U232 ( .A1(n2245), .A2(n2270), .B1(n3146), .B2(n2880), .ZN(n1664)
         );
  OAI22_X1 U233 ( .A1(n2233), .A2(n2270), .B1(n3148), .B2(n2879), .ZN(n1673)
         );
  OAI22_X1 U234 ( .A1(n2248), .A2(n2270), .B1(n3148), .B2(n2869), .ZN(n1663)
         );
  OAI22_X1 U235 ( .A1(n2252), .A2(n2270), .B1(n3146), .B2(n2881), .ZN(n1661)
         );
  OAI22_X1 U236 ( .A1(n2268), .A2(n2270), .B1(n3148), .B2(n2877), .ZN(n1653)
         );
  OAI22_X1 U237 ( .A1(n2210), .A2(n2270), .B1(n3146), .B2(n2863), .ZN(n1684)
         );
  OAI22_X1 U238 ( .A1(n2237), .A2(n2270), .B1(n3149), .B2(n2884), .ZN(n1669)
         );
  OAI22_X1 U239 ( .A1(n2235), .A2(n2270), .B1(n3147), .B2(n2870), .ZN(n1672)
         );
  OAI22_X1 U240 ( .A1(n2231), .A2(n2270), .B1(n3148), .B2(n2883), .ZN(n1674)
         );
  OAI22_X1 U241 ( .A1(n2250), .A2(n2270), .B1(n3146), .B2(n2882), .ZN(n1662)
         );
  OAI22_X1 U243 ( .A1(n2215), .A2(n2270), .B1(n3146), .B2(n2811), .ZN(n1682)
         );
  OAI22_X1 U244 ( .A1(n2266), .A2(n2270), .B1(n3148), .B2(n2878), .ZN(n1654)
         );
  OAI22_X1 U245 ( .A1(n2239), .A2(n2270), .B1(n3147), .B2(n2866), .ZN(n1668)
         );
  OAI22_X1 U246 ( .A1(n2243), .A2(n2270), .B1(n3147), .B2(n2885), .ZN(n1665)
         );
  OAI22_X1 U247 ( .A1(n2229), .A2(n2270), .B1(n3146), .B2(n2871), .ZN(n1675)
         );
  OAI22_X1 U248 ( .A1(n2227), .A2(n2270), .B1(n3148), .B2(n2873), .ZN(n1676)
         );
  OAI22_X1 U249 ( .A1(n2254), .A2(n2270), .B1(n3149), .B2(n2867), .ZN(n1660)
         );
  OAI22_X1 U250 ( .A1(n2225), .A2(n2270), .B1(n3149), .B2(n2800), .ZN(n1677)
         );
  OAI22_X1 U251 ( .A1(n2256), .A2(n2270), .B1(n3147), .B2(n2872), .ZN(n1659)
         );
  OAI22_X1 U252 ( .A1(n2223), .A2(n2270), .B1(n3149), .B2(n2833), .ZN(n1678)
         );
  OAI22_X1 U253 ( .A1(n2221), .A2(n2270), .B1(n3147), .B2(n2822), .ZN(n1679)
         );
  OAI22_X1 U254 ( .A1(n2219), .A2(n2270), .B1(n3149), .B2(n2844), .ZN(n1680)
         );
  OAI22_X1 U255 ( .A1(n2258), .A2(n2270), .B1(n3149), .B2(n2875), .ZN(n1658)
         );
  OAI22_X1 U256 ( .A1(n2260), .A2(n2270), .B1(n3149), .B2(n2874), .ZN(n1657)
         );
  OAI22_X1 U257 ( .A1(n2262), .A2(n2270), .B1(n3148), .B2(n2876), .ZN(n1656)
         );
  OAI22_X1 U258 ( .A1(n2264), .A2(n2270), .B1(n3146), .B2(n2868), .ZN(n1655)
         );
  OAI22_X1 U259 ( .A1(n3151), .A2(n2920), .B1(n2237), .B2(n2994), .ZN(n1701)
         );
  OAI22_X1 U260 ( .A1(n3153), .A2(n2907), .B1(n2239), .B2(n2994), .ZN(n1700)
         );
  OAI22_X1 U261 ( .A1(n3154), .A2(n2921), .B1(n2243), .B2(n2994), .ZN(n1697)
         );
  OAI22_X1 U262 ( .A1(n3150), .A2(n2897), .B1(n2235), .B2(n2994), .ZN(n1704)
         );
  OAI22_X1 U263 ( .A1(n3153), .A2(n2901), .B1(n2245), .B2(n2994), .ZN(n1696)
         );
  OAI22_X1 U264 ( .A1(n3151), .A2(n2906), .B1(n2233), .B2(n2994), .ZN(n1705)
         );
  OAI22_X1 U265 ( .A1(n3152), .A2(n2915), .B1(n2248), .B2(n2994), .ZN(n1695)
         );
  OAI22_X1 U266 ( .A1(n3150), .A2(n2918), .B1(n2250), .B2(n2994), .ZN(n1694)
         );
  OAI22_X1 U267 ( .A1(n3152), .A2(n2916), .B1(n2252), .B2(n2994), .ZN(n1693)
         );
  OAI22_X1 U268 ( .A1(n3152), .A2(n2910), .B1(n2227), .B2(n2993), .ZN(n1708)
         );
  OAI22_X1 U269 ( .A1(n3151), .A2(n2894), .B1(n2254), .B2(n2994), .ZN(n1692)
         );
  OAI22_X1 U270 ( .A1(n3152), .A2(n2902), .B1(n2231), .B2(n2993), .ZN(n1706)
         );
  OAI22_X1 U271 ( .A1(n3154), .A2(n2917), .B1(n2229), .B2(n2994), .ZN(n1707)
         );
  OAI22_X1 U272 ( .A1(n3153), .A2(n2909), .B1(n2225), .B2(n2993), .ZN(n1709)
         );
  OAI22_X1 U273 ( .A1(n3154), .A2(n2895), .B1(n2223), .B2(n2993), .ZN(n1710)
         );
  OAI22_X1 U274 ( .A1(n3150), .A2(n2903), .B1(n2221), .B2(n2993), .ZN(n1711)
         );
  OAI22_X1 U275 ( .A1(n3150), .A2(n2896), .B1(n2219), .B2(n2993), .ZN(n1712)
         );
  OAI22_X1 U276 ( .A1(n3153), .A2(n2904), .B1(n2217), .B2(n2993), .ZN(n1713)
         );
  OAI22_X1 U277 ( .A1(n3151), .A2(n2900), .B1(n2215), .B2(n2993), .ZN(n1714)
         );
  OAI22_X1 U278 ( .A1(n3152), .A2(n2914), .B1(n2213), .B2(n2993), .ZN(n1715)
         );
  OAI22_X1 U279 ( .A1(n3151), .A2(n2913), .B1(n2268), .B2(n2993), .ZN(n1685)
         );
  OAI22_X1 U280 ( .A1(n3150), .A2(n2908), .B1(n2256), .B2(n2995), .ZN(n1691)
         );
  OAI22_X1 U281 ( .A1(n3154), .A2(n2898), .B1(n2258), .B2(n2995), .ZN(n1690)
         );
  OAI22_X1 U282 ( .A1(n3154), .A2(n2911), .B1(n2260), .B2(n2995), .ZN(n1689)
         );
  OAI22_X1 U283 ( .A1(n3151), .A2(n2899), .B1(n2262), .B2(n2995), .ZN(n1688)
         );
  OAI22_X1 U284 ( .A1(n3153), .A2(n2912), .B1(n2264), .B2(n2995), .ZN(n1687)
         );
  OAI22_X1 U285 ( .A1(n3152), .A2(n2905), .B1(n2266), .B2(n2995), .ZN(n1686)
         );
  OAI22_X1 U286 ( .A1(n3153), .A2(n2919), .B1(n2210), .B2(n2994), .ZN(n1716)
         );
  OAI22_X1 U287 ( .A1(n2237), .A2(n2991), .B1(n3142), .B2(n2653), .ZN(n1637)
         );
  OAI22_X1 U288 ( .A1(n2239), .A2(n2991), .B1(n3144), .B2(n2513), .ZN(n1636)
         );
  OAI22_X1 U289 ( .A1(n2223), .A2(n2975), .B1(n3111), .B2(n2888), .ZN(n1454)
         );
  OAI22_X1 U290 ( .A1(n2258), .A2(n2977), .B1(n3112), .B2(n2887), .ZN(n1434)
         );
  OAI22_X1 U291 ( .A1(n2266), .A2(n2977), .B1(n3113), .B2(n2889), .ZN(n1430)
         );
  OAI22_X1 U292 ( .A1(n2215), .A2(n2975), .B1(n3114), .B2(n2890), .ZN(n1458)
         );
  OAI22_X1 U293 ( .A1(n2210), .A2(n2976), .B1(n3114), .B2(n2891), .ZN(n1460)
         );
  OAI22_X1 U294 ( .A1(n2219), .A2(n2990), .B1(n3141), .B2(n2455), .ZN(n1648)
         );
  OAI22_X1 U295 ( .A1(n2235), .A2(n2991), .B1(n3141), .B2(n2457), .ZN(n1640)
         );
  OAI22_X1 U296 ( .A1(n2221), .A2(n2990), .B1(n3141), .B2(n2503), .ZN(n1647)
         );
  OAI22_X1 U297 ( .A1(n2250), .A2(n2991), .B1(n3141), .B2(n2623), .ZN(n1630)
         );
  OAI22_X1 U298 ( .A1(n2256), .A2(n2992), .B1(n3141), .B2(n2514), .ZN(n1627)
         );
  OAI22_X1 U299 ( .A1(n2233), .A2(n2991), .B1(n3142), .B2(n2512), .ZN(n1641)
         );
  OAI22_X1 U300 ( .A1(n2248), .A2(n2991), .B1(n3143), .B2(n2590), .ZN(n1631)
         );
  OAI22_X1 U302 ( .A1(n2254), .A2(n2992), .B1(n3142), .B2(n2450), .ZN(n1628)
         );
  OAI22_X1 U303 ( .A1(n2213), .A2(n2990), .B1(n3143), .B2(n2579), .ZN(n1651)
         );
  OAI22_X1 U304 ( .A1(n2268), .A2(n2990), .B1(n3142), .B2(n2568), .ZN(n1621)
         );
  OAI22_X1 U305 ( .A1(n2252), .A2(n2991), .B1(n3143), .B2(n2601), .ZN(n1629)
         );
  OAI22_X1 U306 ( .A1(n2217), .A2(n2991), .B1(n3144), .B2(n2506), .ZN(n1649)
         );
  OAI22_X1 U307 ( .A1(n2245), .A2(n2991), .B1(n3144), .B2(n2476), .ZN(n1632)
         );
  OAI22_X1 U308 ( .A1(n2231), .A2(n2990), .B1(n3143), .B2(n2498), .ZN(n1642)
         );
  OAI22_X1 U309 ( .A1(n2227), .A2(n2990), .B1(n3143), .B2(n2535), .ZN(n1644)
         );
  OAI22_X1 U310 ( .A1(n2225), .A2(n2990), .B1(n3144), .B2(n2522), .ZN(n1645)
         );
  OAI22_X1 U311 ( .A1(n2215), .A2(n2990), .B1(n3142), .B2(n2472), .ZN(n1650)
         );
  OAI22_X1 U312 ( .A1(n2266), .A2(n2992), .B1(n3143), .B2(n2507), .ZN(n1622)
         );
  OAI22_X1 U313 ( .A1(n2210), .A2(n2991), .B1(n3144), .B2(n2644), .ZN(n1652)
         );
  OAI22_X1 U314 ( .A1(n2264), .A2(n2992), .B1(n3144), .B2(n2557), .ZN(n1623)
         );
  OAI22_X1 U315 ( .A1(n2262), .A2(n2992), .B1(n3142), .B2(n2460), .ZN(n1624)
         );
  OAI22_X1 U316 ( .A1(n2225), .A2(n2975), .B1(n3115), .B2(n2886), .ZN(n1453)
         );
  OAI22_X1 U317 ( .A1(n2229), .A2(n2991), .B1(n3145), .B2(n2612), .ZN(n1643)
         );
  OAI22_X1 U318 ( .A1(n2243), .A2(n2991), .B1(n3145), .B2(n2655), .ZN(n1633)
         );
  OAI22_X1 U319 ( .A1(n2223), .A2(n2990), .B1(n3145), .B2(n2451), .ZN(n1646)
         );
  OAI22_X1 U320 ( .A1(n2258), .A2(n2992), .B1(n3145), .B2(n2458), .ZN(n1626)
         );
  OAI22_X1 U321 ( .A1(n2260), .A2(n2992), .B1(n3145), .B2(n2546), .ZN(n1625)
         );
  INV_X1 U322 ( .A(n2489), .ZN(PRED[15]) );
  AOI222_X1 U323 ( .A1(PRED_TK[15]), .A2(n3091), .B1(NEXT_PC[15]), .B2(n3095), 
        .C1(NEW_PC[15]), .C2(n3101), .ZN(n2489) );
  NAND2_X1 U324 ( .A1(n2666), .A2(n2990), .ZN(n1635) );
  NAND2_X1 U325 ( .A1(n2789), .A2(n2990), .ZN(n1638) );
  NAND2_X1 U326 ( .A1(n2662), .A2(n2990), .ZN(n1634) );
  NAND2_X1 U327 ( .A1(n2892), .A2(n2993), .ZN(n1698) );
  NAND2_X1 U328 ( .A1(n2893), .A2(n2993), .ZN(n1699) );
  BUF_X1 U329 ( .A(INST[15]), .Z(n3182) );
  INV_X1 U330 ( .A(n2493), .ZN(PRED[11]) );
  AOI222_X1 U331 ( .A1(PRED_TK[11]), .A2(n2462), .B1(NEXT_PC[11]), .B2(n3093), 
        .C1(NEW_PC[11]), .C2(n3105), .ZN(n2493) );
  INV_X1 U332 ( .A(n2494), .ZN(PRED[10]) );
  AOI222_X1 U333 ( .A1(PRED_TK[10]), .A2(n3092), .B1(NEXT_PC[10]), .B2(n3095), 
        .C1(NEW_PC[10]), .C2(n3098), .ZN(n2494) );
  INV_X1 U334 ( .A(n2470), .ZN(PRED[3]) );
  AOI222_X1 U335 ( .A1(PRED_TK[3]), .A2(n3092), .B1(NEXT_PC[3]), .B2(n3093), 
        .C1(NEW_PC[3]), .C2(n3098), .ZN(n2470) );
  INV_X1 U336 ( .A(n2469), .ZN(PRED[4]) );
  AOI222_X1 U337 ( .A1(PRED_TK[4]), .A2(n2462), .B1(NEXT_PC[4]), .B2(n3095), 
        .C1(NEW_PC[4]), .C2(n3099), .ZN(n2469) );
  INV_X1 U338 ( .A(n2467), .ZN(PRED[6]) );
  AOI222_X1 U339 ( .A1(PRED_TK[6]), .A2(n3092), .B1(NEXT_PC[6]), .B2(n3095), 
        .C1(NEW_PC[6]), .C2(n3101), .ZN(n2467) );
  INV_X1 U340 ( .A(n2466), .ZN(PRED[7]) );
  AOI222_X1 U341 ( .A1(PRED_TK[7]), .A2(n2462), .B1(NEXT_PC[7]), .B2(n3093), 
        .C1(NEW_PC[7]), .C2(n3096), .ZN(n2466) );
  INV_X1 U342 ( .A(n2490), .ZN(PRED[14]) );
  AOI222_X1 U343 ( .A1(PRED_TK[14]), .A2(n2462), .B1(NEXT_PC[14]), .B2(n3094), 
        .C1(NEW_PC[14]), .C2(n3099), .ZN(n2490) );
  INV_X1 U344 ( .A(n2486), .ZN(PRED[18]) );
  AOI222_X1 U345 ( .A1(PRED_TK[18]), .A2(n3091), .B1(NEXT_PC[18]), .B2(n3094), 
        .C1(NEW_PC[18]), .C2(n3102), .ZN(n2486) );
  INV_X1 U346 ( .A(n2481), .ZN(PRED[22]) );
  AOI222_X1 U347 ( .A1(PRED_TK[22]), .A2(n2462), .B1(NEXT_PC[22]), .B2(n3094), 
        .C1(NEW_PC[22]), .C2(n3096), .ZN(n2481) );
  INV_X1 U348 ( .A(n2477), .ZN(PRED[26]) );
  AOI222_X1 U349 ( .A1(PRED_TK[26]), .A2(n3091), .B1(NEXT_PC[26]), .B2(n3094), 
        .C1(NEW_PC[26]), .C2(n3105), .ZN(n2477) );
  INV_X1 U350 ( .A(n2491), .ZN(PRED[13]) );
  AOI222_X1 U351 ( .A1(PRED_TK[13]), .A2(n3092), .B1(NEXT_PC[13]), .B2(n3094), 
        .C1(NEW_PC[13]), .C2(n3099), .ZN(n2491) );
  INV_X1 U352 ( .A(n2473), .ZN(PRED[2]) );
  AOI222_X1 U353 ( .A1(PRED_TK[2]), .A2(n3092), .B1(NEXT_PC[2]), .B2(n3094), 
        .C1(NEW_PC[2]), .C2(n3104), .ZN(n2473) );
  INV_X1 U354 ( .A(n2468), .ZN(PRED[5]) );
  AOI222_X1 U355 ( .A1(PRED_TK[5]), .A2(n3091), .B1(NEXT_PC[5]), .B2(n3094), 
        .C1(NEW_PC[5]), .C2(n3096), .ZN(n2468) );
  INV_X1 U356 ( .A(n2485), .ZN(PRED[19]) );
  AOI222_X1 U357 ( .A1(PRED_TK[19]), .A2(n3092), .B1(NEXT_PC[19]), .B2(n3095), 
        .C1(NEW_PC[19]), .C2(n3096), .ZN(n2485) );
  INV_X1 U358 ( .A(n2483), .ZN(PRED[20]) );
  AOI222_X1 U359 ( .A1(PRED_TK[20]), .A2(n3091), .B1(NEXT_PC[20]), .B2(n3093), 
        .C1(NEW_PC[20]), .C2(n3104), .ZN(n2483) );
  INV_X1 U360 ( .A(n2480), .ZN(PRED[23]) );
  AOI222_X1 U361 ( .A1(PRED_TK[23]), .A2(n3091), .B1(NEXT_PC[23]), .B2(n3095), 
        .C1(NEW_PC[23]), .C2(n3096), .ZN(n2480) );
  INV_X1 U362 ( .A(n2479), .ZN(PRED[24]) );
  AOI222_X1 U363 ( .A1(PRED_TK[24]), .A2(n3092), .B1(NEXT_PC[24]), .B2(n3093), 
        .C1(NEW_PC[24]), .C2(n3104), .ZN(n2479) );
  INV_X1 U364 ( .A(n2478), .ZN(PRED[25]) );
  AOI222_X1 U366 ( .A1(PRED_TK[25]), .A2(n2462), .B1(NEXT_PC[25]), .B2(n3095), 
        .C1(NEW_PC[25]), .C2(n3104), .ZN(n2478) );
  INV_X1 U367 ( .A(n2475), .ZN(PRED[28]) );
  AOI222_X1 U368 ( .A1(PRED_TK[28]), .A2(n2462), .B1(NEXT_PC[28]), .B2(n3093), 
        .C1(NEW_PC[28]), .C2(n3105), .ZN(n2475) );
  INV_X1 U369 ( .A(n2474), .ZN(PRED[29]) );
  AOI222_X1 U370 ( .A1(PRED_TK[29]), .A2(n3091), .B1(NEXT_PC[29]), .B2(n3093), 
        .C1(NEW_PC[29]), .C2(n3105), .ZN(n2474) );
  INV_X1 U371 ( .A(n2492), .ZN(PRED[12]) );
  AOI222_X1 U372 ( .A1(PRED_TK[12]), .A2(n3091), .B1(NEXT_PC[12]), .B2(n3093), 
        .C1(NEW_PC[12]), .C2(n3099), .ZN(n2492) );
  INV_X1 U373 ( .A(n2488), .ZN(PRED[16]) );
  AOI222_X1 U374 ( .A1(PRED_TK[16]), .A2(n3092), .B1(NEXT_PC[16]), .B2(n3093), 
        .C1(NEW_PC[16]), .C2(n3096), .ZN(n2488) );
  INV_X1 U375 ( .A(n2487), .ZN(PRED[17]) );
  AOI222_X1 U376 ( .A1(PRED_TK[17]), .A2(n2462), .B1(NEXT_PC[17]), .B2(n3095), 
        .C1(NEW_PC[17]), .C2(n3101), .ZN(n2487) );
  INV_X1 U377 ( .A(n2465), .ZN(PRED[8]) );
  AOI222_X1 U378 ( .A1(PRED_TK[8]), .A2(n3091), .B1(NEXT_PC[8]), .B2(n3093), 
        .C1(NEW_PC[8]), .C2(n3096), .ZN(n2465) );
  OAI221_X1 U379 ( .B1(n2496), .B2(n2497), .C1(n2362), .C2(n2407), .A(n2114), 
        .ZN(n2463) );
  NAND3_X1 U380 ( .A1(n2996), .A2(n2997), .A3(n2998), .ZN(PRED[30]) );
  NOR2_X1 U381 ( .A1(n2860), .A2(n2855), .ZN(n2849) );
  NOR2_X1 U382 ( .A1(n2861), .A2(n2862), .ZN(n2847) );
  NAND2_X1 U383 ( .A1(n2853), .A2(n2854), .ZN(n3018) );
  NAND2_X1 U384 ( .A1(n2853), .A2(n2854), .ZN(n3017) );
  NAND2_X1 U385 ( .A1(n2853), .A2(n2850), .ZN(n3083) );
  NAND2_X1 U386 ( .A1(n2846), .A2(n2847), .ZN(n2332) );
  NAND2_X1 U387 ( .A1(n2846), .A2(n2847), .ZN(n3090) );
  NAND2_X1 U388 ( .A1(n2846), .A2(n2848), .ZN(n3088) );
  NAND2_X1 U389 ( .A1(n2846), .A2(n2847), .ZN(n3089) );
  NAND2_X1 U390 ( .A1(n2846), .A2(n2848), .ZN(n3087) );
  NAND2_X1 U391 ( .A1(n2853), .A2(n2854), .ZN(n2349) );
  NAND2_X1 U392 ( .A1(n2853), .A2(n2850), .ZN(n3084) );
  NAND2_X1 U393 ( .A1(n2853), .A2(n2850), .ZN(n2343) );
  NAND2_X1 U394 ( .A1(n2846), .A2(n2848), .ZN(n2269) );
  AND2_X1 U395 ( .A1(n2850), .A2(n2851), .ZN(n2081) );
  AND2_X1 U396 ( .A1(n2850), .A2(n2851), .ZN(n3086) );
  AND2_X1 U397 ( .A1(n2850), .A2(n2851), .ZN(n3085) );
  OAI22_X1 U398 ( .A1(n2269), .A2(n2894), .B1(n2332), .B2(n2450), .ZN(n2790)
         );
  OAI22_X1 U399 ( .A1(n2269), .A2(n2895), .B1(n2332), .B2(n2451), .ZN(n2823)
         );
  OAI22_X1 U400 ( .A1(n3088), .A2(n2896), .B1(n2332), .B2(n2455), .ZN(n2536)
         );
  OAI22_X1 U401 ( .A1(n2269), .A2(n2897), .B1(n2332), .B2(n2457), .ZN(n2691)
         );
  OAI22_X1 U402 ( .A1(n3088), .A2(n2898), .B1(n3090), .B2(n2458), .ZN(n2834)
         );
  OAI22_X1 U403 ( .A1(n3087), .A2(n2899), .B1(n3090), .B2(n2460), .ZN(n2547)
         );
  OAI22_X1 U404 ( .A1(n3087), .A2(n2900), .B1(n3090), .B2(n2472), .ZN(n2580)
         );
  OAI22_X1 U405 ( .A1(n3088), .A2(n2901), .B1(n3090), .B2(n2476), .ZN(n2702)
         );
  OAI22_X1 U406 ( .A1(n3088), .A2(n2902), .B1(n3090), .B2(n2498), .ZN(n2735)
         );
  OAI22_X1 U407 ( .A1(n3088), .A2(n2892), .B1(n3090), .B2(n2662), .ZN(n2667)
         );
  OAI22_X1 U408 ( .A1(n3087), .A2(n2903), .B1(n3089), .B2(n2503), .ZN(n2845)
         );
  OAI22_X1 U409 ( .A1(n2269), .A2(n2904), .B1(n3089), .B2(n2506), .ZN(n2558)
         );
  OAI22_X1 U410 ( .A1(n2269), .A2(n2905), .B1(n3089), .B2(n2507), .ZN(n2591)
         );
  OAI22_X1 U411 ( .A1(n3087), .A2(n2906), .B1(n3089), .B2(n2512), .ZN(n2713)
         );
  OAI22_X1 U412 ( .A1(n2269), .A2(n2893), .B1(n3089), .B2(n2666), .ZN(n2654)
         );
  OAI22_X1 U413 ( .A1(n3079), .A2(n2800), .B1(n3083), .B2(n2668), .ZN(n2802)
         );
  OAI22_X1 U414 ( .A1(n3080), .A2(n2811), .B1(n3083), .B2(n2679), .ZN(n2581)
         );
  OAI22_X1 U415 ( .A1(n3081), .A2(n2822), .B1(n3084), .B2(n2690), .ZN(n2852)
         );
  OAI22_X1 U416 ( .A1(n3079), .A2(n2833), .B1(n2343), .B2(n2701), .ZN(n2824)
         );
  OAI22_X1 U417 ( .A1(n3081), .A2(n2844), .B1(n2343), .B2(n2712), .ZN(n2537)
         );
  OAI22_X1 U418 ( .A1(n3079), .A2(n2863), .B1(n3084), .B2(n2723), .ZN(n2625)
         );
  NAND2_X1 U419 ( .A1(n2846), .A2(n2854), .ZN(n2298) );
  NAND4_X1 U420 ( .A1(n2499), .A2(n2500), .A3(n2501), .A4(n2502), .ZN(n2497)
         );
  AOI221_X1 U421 ( .B1(n2509), .B2(n2948), .C1(n2510), .C2(n2745), .A(n2511), 
        .ZN(n2500) );
  AOI221_X1 U422 ( .B1(n3000), .B2(n2412), .C1(n3009), .C2(n2447), .A(n2515), 
        .ZN(n2499) );
  AOI221_X1 U423 ( .B1(n3051), .B2(n2951), .C1(n3076), .C2(n2767), .A(n2508), 
        .ZN(n2501) );
  NAND2_X1 U424 ( .A1(n2853), .A2(n2848), .ZN(n2346) );
  NAND2_X1 U425 ( .A1(n2853), .A2(n2847), .ZN(n2352) );
  NAND2_X1 U426 ( .A1(n2850), .A2(n2849), .ZN(n2355) );
  NAND2_X1 U427 ( .A1(n2850), .A2(n2849), .ZN(n3033) );
  NAND2_X1 U428 ( .A1(n2848), .A2(n2851), .ZN(n2113) );
  NAND2_X1 U430 ( .A1(n2854), .A2(n2849), .ZN(n3019) );
  NAND2_X1 U431 ( .A1(n2854), .A2(n2849), .ZN(n2371) );
  NAND2_X1 U432 ( .A1(n2848), .A2(n2849), .ZN(n2368) );
  NAND2_X1 U433 ( .A1(n2848), .A2(n2849), .ZN(n3026) );
  NAND2_X1 U434 ( .A1(n2851), .A2(n2847), .ZN(n2176) );
  AND2_X1 U435 ( .A1(n2854), .A2(n2851), .ZN(n2145) );
  AND2_X1 U436 ( .A1(n2854), .A2(n2851), .ZN(n3063) );
  AND2_X1 U437 ( .A1(n2846), .A2(n2850), .ZN(n3050) );
  AND2_X1 U438 ( .A1(n2846), .A2(n2850), .ZN(n2207) );
  AND2_X1 U439 ( .A1(n2846), .A2(n2850), .ZN(n3049) );
  NAND2_X1 U440 ( .A1(n2423), .A2(n2420), .ZN(n2375) );
  NAND2_X1 U441 ( .A1(n2422), .A2(n2416), .ZN(n2405) );
  NAND2_X1 U442 ( .A1(n2422), .A2(n2418), .ZN(n2401) );
  NAND2_X1 U443 ( .A1(n2422), .A2(n2419), .ZN(n2397) );
  NAND2_X1 U444 ( .A1(n2422), .A2(n2420), .ZN(n2393) );
  NAND2_X1 U445 ( .A1(n2417), .A2(n2420), .ZN(n2391) );
  NAND2_X1 U446 ( .A1(n2415), .A2(n2420), .ZN(n2389) );
  NAND2_X1 U447 ( .A1(n2417), .A2(n2419), .ZN(n2387) );
  NAND2_X1 U448 ( .A1(n2415), .A2(n2419), .ZN(n2385) );
  NAND2_X1 U449 ( .A1(n2417), .A2(n2418), .ZN(n2383) );
  NAND2_X1 U450 ( .A1(n2415), .A2(n2418), .ZN(n2381) );
  NAND2_X1 U451 ( .A1(n2417), .A2(n2416), .ZN(n2379) );
  NAND2_X1 U452 ( .A1(n2415), .A2(n2416), .ZN(n2377) );
  INV_X1 U453 ( .A(n2424), .ZN(n2418) );
  INV_X1 U454 ( .A(n2425), .ZN(n2416) );
  NAND2_X1 U455 ( .A1(n2419), .A2(n2423), .ZN(n2395) );
  NAND2_X1 U456 ( .A1(n2416), .A2(n2423), .ZN(n2403) );
  NAND2_X1 U457 ( .A1(n2418), .A2(n2423), .ZN(n2399) );
  INV_X1 U458 ( .A(n2419), .ZN(n2449) );
  OAI22_X2 U459 ( .A1(n2406), .A2(n2407), .B1(n2408), .B2(n2426), .ZN(n2414)
         );
  AOI22_X1 U460 ( .A1(n2411), .A2(n2421), .B1(n747), .B2(n2413), .ZN(n2426) );
  OAI22_X2 U461 ( .A1(n2406), .A2(n2407), .B1(n2408), .B2(n2409), .ZN(n2374)
         );
  INV_X1 U462 ( .A(n2410), .ZN(n2409) );
  OAI22_X1 U463 ( .A1(n2411), .A2(n747), .B1(n2421), .B2(n2413), .ZN(n2410) );
  INV_X1 U464 ( .A(n2495), .ZN(PRED[0]) );
  AOI222_X1 U465 ( .A1(PRED_TK[0]), .A2(n3091), .B1(NEXT_PC[0]), .B2(n3094), 
        .C1(NEW_PC[0]), .C2(n3104), .ZN(n2495) );
  OAI22_X1 U466 ( .A1(n992), .A2(n3138), .B1(n2237), .B2(n2335), .ZN(n1605) );
  OAI22_X1 U467 ( .A1(n988), .A2(n3137), .B1(n2243), .B2(n2335), .ZN(n1601) );
  OAI22_X1 U468 ( .A1(n995), .A2(n3138), .B1(n2235), .B2(n2335), .ZN(n1608) );
  OAI22_X1 U469 ( .A1(n987), .A2(n3136), .B1(n2245), .B2(n2335), .ZN(n1600) );
  OAI22_X1 U470 ( .A1(n996), .A2(n3139), .B1(n2233), .B2(n2335), .ZN(n1609) );
  OAI22_X1 U471 ( .A1(n986), .A2(n3137), .B1(n2248), .B2(n2335), .ZN(n1599) );
  OAI22_X1 U472 ( .A1(n985), .A2(n3137), .B1(n2250), .B2(n2335), .ZN(n1598) );
  OAI22_X1 U473 ( .A1(n998), .A2(n3136), .B1(n2229), .B2(n2335), .ZN(n1611) );
  OAI22_X1 U474 ( .A1(n984), .A2(n3140), .B1(n2252), .B2(n2335), .ZN(n1597) );
  OAI22_X1 U475 ( .A1(n991), .A2(n3138), .B1(n2239), .B2(n2335), .ZN(n1604) );
  OAI22_X1 U476 ( .A1(n997), .A2(n3140), .B1(n2231), .B2(n2335), .ZN(n1610) );
  OAI22_X1 U477 ( .A1(n999), .A2(n3139), .B1(n2227), .B2(n2335), .ZN(n1612) );
  OAI22_X1 U478 ( .A1(n976), .A2(n3140), .B1(n2268), .B2(n2335), .ZN(n1589) );
  OAI22_X1 U479 ( .A1(n983), .A2(n3139), .B1(n2254), .B2(n2335), .ZN(n1596) );
  OAI22_X1 U480 ( .A1(n982), .A2(n3138), .B1(n2256), .B2(n2335), .ZN(n1595) );
  OAI22_X1 U481 ( .A1(n981), .A2(n3136), .B1(n2258), .B2(n2335), .ZN(n1594) );
  OAI22_X1 U482 ( .A1(n980), .A2(n3136), .B1(n2260), .B2(n2335), .ZN(n1593) );
  OAI22_X1 U483 ( .A1(n979), .A2(n3137), .B1(n2262), .B2(n2335), .ZN(n1592) );
  OAI22_X1 U484 ( .A1(n978), .A2(n3136), .B1(n2264), .B2(n2335), .ZN(n1591) );
  OAI22_X1 U485 ( .A1(n977), .A2(n3140), .B1(n2266), .B2(n2335), .ZN(n1590) );
  OAI22_X1 U486 ( .A1(n2217), .A2(n2270), .B1(n1068), .B2(n3147), .ZN(n1681)
         );
  OAI22_X1 U487 ( .A1(n2213), .A2(n2270), .B1(n1070), .B2(n3146), .ZN(n1683)
         );
  OAI22_X1 U488 ( .A1(n960), .A2(n3131), .B1(n2237), .B2(n2988), .ZN(n1573) );
  OAI22_X1 U489 ( .A1(n959), .A2(n3132), .B1(n2239), .B2(n2988), .ZN(n1572) );
  OAI22_X1 U490 ( .A1(n746), .A2(n2376), .B1(n2374), .B2(n2377), .ZN(n1295) );
  OAI22_X1 U491 ( .A1(n732), .A2(n2404), .B1(n2374), .B2(n2405), .ZN(n1281) );
  OAI22_X1 U492 ( .A1(n745), .A2(n2378), .B1(n2374), .B2(n2379), .ZN(n1294) );
  OAI22_X1 U493 ( .A1(n733), .A2(n2402), .B1(n2374), .B2(n2403), .ZN(n1282) );
  OAI22_X1 U494 ( .A1(n744), .A2(n2380), .B1(n2374), .B2(n2381), .ZN(n1293) );
  OAI22_X1 U495 ( .A1(n734), .A2(n2400), .B1(n2374), .B2(n2401), .ZN(n1283) );
  OAI22_X1 U496 ( .A1(n743), .A2(n2382), .B1(n2374), .B2(n2383), .ZN(n1292) );
  OAI22_X1 U497 ( .A1(n735), .A2(n2398), .B1(n2374), .B2(n2399), .ZN(n1284) );
  OAI22_X1 U498 ( .A1(n742), .A2(n2384), .B1(n2374), .B2(n2385), .ZN(n1291) );
  OAI22_X1 U499 ( .A1(n736), .A2(n2396), .B1(n2374), .B2(n2397), .ZN(n1285) );
  OAI22_X1 U500 ( .A1(n741), .A2(n2386), .B1(n2374), .B2(n2387), .ZN(n1290) );
  OAI22_X1 U501 ( .A1(n737), .A2(n2394), .B1(n2374), .B2(n2395), .ZN(n1286) );
  OAI22_X1 U502 ( .A1(n740), .A2(n2388), .B1(n2374), .B2(n2389), .ZN(n1289) );
  OAI22_X1 U503 ( .A1(n738), .A2(n2392), .B1(n2374), .B2(n2393), .ZN(n1287) );
  OAI22_X1 U504 ( .A1(n739), .A2(n2390), .B1(n2374), .B2(n2391), .ZN(n1288) );
  OAI22_X1 U505 ( .A1(n752), .A2(n2373), .B1(n2374), .B2(n2375), .ZN(n1360) );
  OAI22_X1 U506 ( .A1(n956), .A2(n3134), .B1(n2243), .B2(n2988), .ZN(n1569) );
  OAI22_X1 U507 ( .A1(n963), .A2(n3135), .B1(n2235), .B2(n2988), .ZN(n1576) );
  OAI22_X1 U508 ( .A1(n955), .A2(n3133), .B1(n2245), .B2(n2988), .ZN(n1568) );
  OAI22_X1 U509 ( .A1(n964), .A2(n3131), .B1(n2233), .B2(n2988), .ZN(n1577) );
  OAI22_X1 U510 ( .A1(n954), .A2(n3132), .B1(n2248), .B2(n2988), .ZN(n1567) );
  OAI22_X1 U511 ( .A1(n953), .A2(n3135), .B1(n2250), .B2(n2988), .ZN(n1566) );
  OAI22_X1 U512 ( .A1(n952), .A2(n3131), .B1(n2252), .B2(n2988), .ZN(n1565) );
  OAI22_X1 U513 ( .A1(n967), .A2(n3132), .B1(n2227), .B2(n2988), .ZN(n1580) );
  OAI22_X1 U514 ( .A1(n951), .A2(n3131), .B1(n2254), .B2(n2988), .ZN(n1564) );
  OAI22_X1 U515 ( .A1(n965), .A2(n3132), .B1(n2231), .B2(n2987), .ZN(n1578) );
  OAI22_X1 U516 ( .A1(n966), .A2(n3133), .B1(n2229), .B2(n2987), .ZN(n1579) );
  OAI22_X1 U517 ( .A1(n968), .A2(n3133), .B1(n2225), .B2(n2987), .ZN(n1581) );
  OAI22_X1 U518 ( .A1(n969), .A2(n3134), .B1(n2223), .B2(n2987), .ZN(n1582) );
  OAI22_X1 U519 ( .A1(n970), .A2(n3135), .B1(n2221), .B2(n2987), .ZN(n1583) );
  OAI22_X1 U520 ( .A1(n971), .A2(n3134), .B1(n2219), .B2(n2987), .ZN(n1584) );
  OAI22_X1 U521 ( .A1(n972), .A2(n3133), .B1(n2217), .B2(n2987), .ZN(n1585) );
  OAI22_X1 U522 ( .A1(n973), .A2(n3131), .B1(n2215), .B2(n2987), .ZN(n1586) );
  OAI22_X1 U523 ( .A1(n974), .A2(n3132), .B1(n2213), .B2(n2987), .ZN(n1587) );
  OAI22_X1 U524 ( .A1(n944), .A2(n3131), .B1(n2268), .B2(n2987), .ZN(n1557) );
  OAI22_X1 U525 ( .A1(n950), .A2(n3135), .B1(n2256), .B2(n2989), .ZN(n1563) );
  OAI22_X1 U526 ( .A1(n949), .A2(n3134), .B1(n2258), .B2(n2989), .ZN(n1562) );
  OAI22_X1 U527 ( .A1(n948), .A2(n3134), .B1(n2260), .B2(n2989), .ZN(n1561) );
  OAI22_X1 U528 ( .A1(n947), .A2(n3135), .B1(n2262), .B2(n2989), .ZN(n1560) );
  OAI22_X1 U529 ( .A1(n946), .A2(n3133), .B1(n2264), .B2(n2989), .ZN(n1559) );
  OAI22_X1 U530 ( .A1(n945), .A2(n3132), .B1(n2266), .B2(n2989), .ZN(n1558) );
  OAI22_X1 U531 ( .A1(n975), .A2(n3133), .B1(n2210), .B2(n2988), .ZN(n1588) );
  OAI22_X1 U532 ( .A1(n716), .A2(n2373), .B1(n2375), .B2(n2414), .ZN(n1265) );
  OAI22_X1 U533 ( .A1(n717), .A2(n2404), .B1(n2405), .B2(n2414), .ZN(n1266) );
  OAI22_X1 U534 ( .A1(n718), .A2(n2402), .B1(n2403), .B2(n2414), .ZN(n1267) );
  OAI22_X1 U535 ( .A1(n719), .A2(n2400), .B1(n2401), .B2(n2414), .ZN(n1268) );
  OAI22_X1 U536 ( .A1(n720), .A2(n2398), .B1(n2399), .B2(n2414), .ZN(n1269) );
  OAI22_X1 U537 ( .A1(n721), .A2(n2396), .B1(n2397), .B2(n2414), .ZN(n1270) );
  OAI22_X1 U538 ( .A1(n722), .A2(n2394), .B1(n2395), .B2(n2414), .ZN(n1271) );
  OAI22_X1 U539 ( .A1(n723), .A2(n2392), .B1(n2393), .B2(n2414), .ZN(n1272) );
  OAI22_X1 U540 ( .A1(n724), .A2(n2390), .B1(n2391), .B2(n2414), .ZN(n1273) );
  OAI22_X1 U541 ( .A1(n725), .A2(n2388), .B1(n2389), .B2(n2414), .ZN(n1274) );
  OAI22_X1 U542 ( .A1(n726), .A2(n2386), .B1(n2387), .B2(n2414), .ZN(n1275) );
  OAI22_X1 U543 ( .A1(n727), .A2(n2384), .B1(n2385), .B2(n2414), .ZN(n1276) );
  OAI22_X1 U544 ( .A1(n728), .A2(n2382), .B1(n2383), .B2(n2414), .ZN(n1277) );
  OAI22_X1 U545 ( .A1(n729), .A2(n2380), .B1(n2381), .B2(n2414), .ZN(n1278) );
  OAI22_X1 U546 ( .A1(n730), .A2(n2378), .B1(n2379), .B2(n2414), .ZN(n1279) );
  OAI22_X1 U547 ( .A1(n731), .A2(n2376), .B1(n2377), .B2(n2414), .ZN(n1280) );
  OAI22_X1 U548 ( .A1(n2237), .A2(n2973), .B1(n800), .B2(n3106), .ZN(n1413) );
  OAI22_X1 U549 ( .A1(n2237), .A2(n2982), .B1(n896), .B2(n3121), .ZN(n1509) );
  OAI22_X1 U550 ( .A1(n2237), .A2(n2979), .B1(n864), .B2(n3116), .ZN(n1477) );
  OAI22_X1 U551 ( .A1(n2237), .A2(n2976), .B1(n832), .B2(n3112), .ZN(n1445) );
  OAI22_X1 U552 ( .A1(n2237), .A2(n2985), .B1(n928), .B2(n3126), .ZN(n1541) );
  OAI22_X1 U553 ( .A1(n2239), .A2(n2973), .B1(n799), .B2(n3107), .ZN(n1412) );
  OAI22_X1 U554 ( .A1(n2239), .A2(n2982), .B1(n895), .B2(n3122), .ZN(n1508) );
  OAI22_X1 U555 ( .A1(n2239), .A2(n2979), .B1(n863), .B2(n3117), .ZN(n1476) );
  OAI22_X1 U556 ( .A1(n2239), .A2(n2976), .B1(n831), .B2(n3111), .ZN(n1444) );
  OAI22_X1 U557 ( .A1(n2239), .A2(n2985), .B1(n927), .B2(n3127), .ZN(n1540) );
  OAI22_X1 U558 ( .A1(n2245), .A2(n2973), .B1(n795), .B2(n3108), .ZN(n1408) );
  OAI22_X1 U559 ( .A1(n2233), .A2(n2973), .B1(n804), .B2(n3106), .ZN(n1417) );
  OAI22_X1 U560 ( .A1(n2248), .A2(n2973), .B1(n794), .B2(n3107), .ZN(n1407) );
  OAI22_X1 U561 ( .A1(n2231), .A2(n2972), .B1(n805), .B2(n3107), .ZN(n1418) );
  OAI22_X1 U562 ( .A1(n2229), .A2(n2973), .B1(n806), .B2(n3108), .ZN(n1419) );
  OAI22_X1 U563 ( .A1(n2252), .A2(n2973), .B1(n792), .B2(n3106), .ZN(n1405) );
  OAI22_X1 U564 ( .A1(n2227), .A2(n2972), .B1(n807), .B2(n3107), .ZN(n1420) );
  OAI22_X1 U565 ( .A1(n2254), .A2(n2974), .B1(n791), .B2(n3106), .ZN(n1404) );
  OAI22_X1 U566 ( .A1(n2225), .A2(n2972), .B1(n808), .B2(n3108), .ZN(n1421) );
  OAI22_X1 U567 ( .A1(n2217), .A2(n2973), .B1(n812), .B2(n3108), .ZN(n1425) );
  OAI22_X1 U568 ( .A1(n2215), .A2(n2972), .B1(n813), .B2(n3106), .ZN(n1426) );
  OAI22_X1 U569 ( .A1(n2266), .A2(n2974), .B1(n785), .B2(n3107), .ZN(n1398) );
  OAI22_X1 U570 ( .A1(n2213), .A2(n2972), .B1(n814), .B2(n3107), .ZN(n1427) );
  OAI22_X1 U571 ( .A1(n2268), .A2(n2972), .B1(n784), .B2(n3106), .ZN(n1397) );
  OAI22_X1 U572 ( .A1(n2210), .A2(n2973), .B1(n815), .B2(n3108), .ZN(n1428) );
  OAI22_X1 U573 ( .A1(n2264), .A2(n2974), .B1(n786), .B2(n3108), .ZN(n1399) );
  OAI22_X1 U574 ( .A1(n2233), .A2(n2982), .B1(n900), .B2(n3121), .ZN(n1513) );
  OAI22_X1 U575 ( .A1(n2248), .A2(n2982), .B1(n890), .B2(n3122), .ZN(n1503) );
  OAI22_X1 U576 ( .A1(n2229), .A2(n2982), .B1(n902), .B2(n3123), .ZN(n1515) );
  OAI22_X1 U577 ( .A1(n2254), .A2(n2983), .B1(n887), .B2(n3121), .ZN(n1500) );
  OAI22_X1 U578 ( .A1(n2213), .A2(n2981), .B1(n910), .B2(n3122), .ZN(n1523) );
  OAI22_X1 U579 ( .A1(n2268), .A2(n2981), .B1(n880), .B2(n3121), .ZN(n1493) );
  OAI22_X1 U580 ( .A1(n2245), .A2(n2979), .B1(n859), .B2(n3118), .ZN(n1472) );
  OAI22_X1 U581 ( .A1(n2233), .A2(n2979), .B1(n868), .B2(n3116), .ZN(n1481) );
  OAI22_X1 U582 ( .A1(n2248), .A2(n2979), .B1(n858), .B2(n3117), .ZN(n1471) );
  OAI22_X1 U583 ( .A1(n2252), .A2(n2979), .B1(n856), .B2(n3116), .ZN(n1469) );
  OAI22_X1 U584 ( .A1(n2217), .A2(n2978), .B1(n876), .B2(n3118), .ZN(n1489) );
  OAI22_X1 U585 ( .A1(n2213), .A2(n2978), .B1(n878), .B2(n3117), .ZN(n1491) );
  OAI22_X1 U586 ( .A1(n2268), .A2(n2978), .B1(n848), .B2(n3116), .ZN(n1461) );
  OAI22_X1 U587 ( .A1(n2210), .A2(n2979), .B1(n879), .B2(n3118), .ZN(n1492) );
  OAI22_X1 U588 ( .A1(n2252), .A2(n2982), .B1(n888), .B2(n3121), .ZN(n1501) );
  OAI22_X1 U589 ( .A1(n2217), .A2(n2982), .B1(n908), .B2(n3123), .ZN(n1521) );
  OAI22_X1 U590 ( .A1(n2245), .A2(n2982), .B1(n891), .B2(n3123), .ZN(n1504) );
  OAI22_X1 U591 ( .A1(n2231), .A2(n2981), .B1(n901), .B2(n3122), .ZN(n1514) );
  OAI22_X1 U592 ( .A1(n2227), .A2(n2981), .B1(n903), .B2(n3122), .ZN(n1516) );
  OAI22_X1 U593 ( .A1(n2225), .A2(n2981), .B1(n904), .B2(n3123), .ZN(n1517) );
  OAI22_X1 U594 ( .A1(n2215), .A2(n2981), .B1(n909), .B2(n3121), .ZN(n1522) );
  OAI22_X1 U595 ( .A1(n2266), .A2(n2983), .B1(n881), .B2(n3122), .ZN(n1494) );
  OAI22_X1 U596 ( .A1(n2210), .A2(n2982), .B1(n911), .B2(n3123), .ZN(n1524) );
  OAI22_X1 U597 ( .A1(n2231), .A2(n2978), .B1(n869), .B2(n3117), .ZN(n1482) );
  OAI22_X1 U598 ( .A1(n2215), .A2(n2978), .B1(n877), .B2(n3116), .ZN(n1490) );
  OAI22_X1 U599 ( .A1(n2266), .A2(n2980), .B1(n849), .B2(n3117), .ZN(n1462) );
  OAI22_X1 U600 ( .A1(n2229), .A2(n2978), .B1(n870), .B2(n3118), .ZN(n1483) );
  OAI22_X1 U601 ( .A1(n2227), .A2(n2979), .B1(n871), .B2(n3117), .ZN(n1484) );
  OAI22_X1 U602 ( .A1(n2254), .A2(n2979), .B1(n855), .B2(n3116), .ZN(n1468) );
  OAI22_X1 U603 ( .A1(n2225), .A2(n2978), .B1(n872), .B2(n3118), .ZN(n1485) );
  OAI22_X1 U604 ( .A1(n2245), .A2(n2985), .B1(n923), .B2(n3128), .ZN(n1536) );
  OAI22_X1 U605 ( .A1(n2233), .A2(n2985), .B1(n932), .B2(n3126), .ZN(n1545) );
  OAI22_X1 U606 ( .A1(n2248), .A2(n2985), .B1(n922), .B2(n3127), .ZN(n1535) );
  OAI22_X1 U607 ( .A1(n2252), .A2(n2985), .B1(n920), .B2(n3126), .ZN(n1533) );
  OAI22_X1 U608 ( .A1(n2217), .A2(n2984), .B1(n940), .B2(n3128), .ZN(n1553) );
  OAI22_X1 U609 ( .A1(n2213), .A2(n2984), .B1(n942), .B2(n3127), .ZN(n1555) );
  OAI22_X1 U610 ( .A1(n2268), .A2(n2984), .B1(n912), .B2(n3126), .ZN(n1525) );
  OAI22_X1 U611 ( .A1(n2210), .A2(n2985), .B1(n943), .B2(n3128), .ZN(n1556) );
  OAI22_X1 U612 ( .A1(n2231), .A2(n2984), .B1(n933), .B2(n3127), .ZN(n1546) );
  OAI22_X1 U613 ( .A1(n2215), .A2(n2984), .B1(n941), .B2(n3126), .ZN(n1554) );
  OAI22_X1 U614 ( .A1(n2229), .A2(n2984), .B1(n934), .B2(n3128), .ZN(n1547) );
  OAI22_X1 U615 ( .A1(n2227), .A2(n2985), .B1(n935), .B2(n3127), .ZN(n1548) );
  OAI22_X1 U616 ( .A1(n2254), .A2(n2985), .B1(n919), .B2(n3126), .ZN(n1532) );
  OAI22_X1 U617 ( .A1(n2225), .A2(n2984), .B1(n936), .B2(n3128), .ZN(n1549) );
  OAI22_X1 U618 ( .A1(n2264), .A2(n2983), .B1(n882), .B2(n3123), .ZN(n1495) );
  OAI22_X1 U619 ( .A1(n2264), .A2(n2980), .B1(n850), .B2(n3118), .ZN(n1463) );
  OAI22_X1 U620 ( .A1(n2266), .A2(n2986), .B1(n913), .B2(n3127), .ZN(n1526) );
  OAI22_X1 U621 ( .A1(n2264), .A2(n2986), .B1(n914), .B2(n3128), .ZN(n1527) );
  OAI22_X1 U622 ( .A1(n2243), .A2(n2973), .B1(n796), .B2(n3109), .ZN(n1409) );
  OAI22_X1 U623 ( .A1(n2223), .A2(n2972), .B1(n809), .B2(n3109), .ZN(n1422) );
  OAI22_X1 U624 ( .A1(n2260), .A2(n2974), .B1(n788), .B2(n3109), .ZN(n1401) );
  OAI22_X1 U625 ( .A1(n2219), .A2(n2972), .B1(n811), .B2(n3109), .ZN(n1424) );
  OAI22_X1 U626 ( .A1(n2258), .A2(n2974), .B1(n789), .B2(n3109), .ZN(n1402) );
  OAI22_X1 U627 ( .A1(n2219), .A2(n2981), .B1(n907), .B2(n3124), .ZN(n1520) );
  OAI22_X1 U628 ( .A1(n2243), .A2(n2982), .B1(n892), .B2(n3124), .ZN(n1505) );
  OAI22_X1 U629 ( .A1(n2223), .A2(n2981), .B1(n905), .B2(n3124), .ZN(n1518) );
  OAI22_X1 U630 ( .A1(n2260), .A2(n2983), .B1(n884), .B2(n3124), .ZN(n1497) );
  OAI22_X1 U631 ( .A1(n2243), .A2(n2979), .B1(n860), .B2(n3119), .ZN(n1473) );
  OAI22_X1 U632 ( .A1(n2223), .A2(n2978), .B1(n873), .B2(n3119), .ZN(n1486) );
  OAI22_X1 U633 ( .A1(n2219), .A2(n2978), .B1(n875), .B2(n3119), .ZN(n1488) );
  OAI22_X1 U634 ( .A1(n2243), .A2(n2985), .B1(n924), .B2(n3129), .ZN(n1537) );
  OAI22_X1 U635 ( .A1(n2223), .A2(n2984), .B1(n937), .B2(n3129), .ZN(n1550) );
  OAI22_X1 U636 ( .A1(n2258), .A2(n2986), .B1(n917), .B2(n3129), .ZN(n1530) );
  OAI22_X1 U637 ( .A1(n2219), .A2(n2984), .B1(n939), .B2(n3129), .ZN(n1552) );
  OAI22_X1 U638 ( .A1(n2258), .A2(n2983), .B1(n885), .B2(n3124), .ZN(n1498) );
  OAI22_X1 U639 ( .A1(n2258), .A2(n2980), .B1(n853), .B2(n3119), .ZN(n1466) );
  OAI22_X1 U640 ( .A1(n2260), .A2(n2980), .B1(n852), .B2(n3119), .ZN(n1465) );
  OAI22_X1 U641 ( .A1(n2260), .A2(n2986), .B1(n916), .B2(n3129), .ZN(n1529) );
  OAI22_X1 U642 ( .A1(n2233), .A2(n2976), .B1(n836), .B2(n3113), .ZN(n1449) );
  OAI22_X1 U643 ( .A1(n2248), .A2(n2976), .B1(n826), .B2(n3111), .ZN(n1439) );
  OAI22_X1 U644 ( .A1(n2229), .A2(n2976), .B1(n838), .B2(n3113), .ZN(n1451) );
  OAI22_X1 U645 ( .A1(n2254), .A2(n2977), .B1(n823), .B2(n3113), .ZN(n1436) );
  OAI22_X1 U646 ( .A1(n2268), .A2(n2975), .B1(n816), .B2(n3111), .ZN(n1429) );
  OAI22_X1 U647 ( .A1(n2235), .A2(n2976), .B1(n835), .B2(n3112), .ZN(n1448) );
  OAI22_X1 U648 ( .A1(n2221), .A2(n2975), .B1(n842), .B2(n3113), .ZN(n1455) );
  OAI22_X1 U649 ( .A1(n2245), .A2(n2976), .B1(n827), .B2(n3112), .ZN(n1440) );
  OAI22_X1 U650 ( .A1(n2231), .A2(n2975), .B1(n837), .B2(n3112), .ZN(n1450) );
  OAI22_X1 U651 ( .A1(n2250), .A2(n2976), .B1(n825), .B2(n3111), .ZN(n1438) );
  OAI22_X1 U652 ( .A1(n2227), .A2(n2975), .B1(n839), .B2(n3113), .ZN(n1452) );
  OAI22_X1 U653 ( .A1(n2264), .A2(n2977), .B1(n818), .B2(n3112), .ZN(n1431) );
  OAI22_X1 U654 ( .A1(n2256), .A2(n2977), .B1(n822), .B2(n3111), .ZN(n1435) );
  OAI22_X1 U655 ( .A1(n2219), .A2(n2975), .B1(n843), .B2(n3114), .ZN(n1456) );
  OAI22_X1 U656 ( .A1(n2252), .A2(n2976), .B1(n824), .B2(n3114), .ZN(n1437) );
  OAI22_X1 U657 ( .A1(n2217), .A2(n2976), .B1(n844), .B2(n3114), .ZN(n1457) );
  OAI22_X1 U658 ( .A1(n3173), .A2(n2237), .B1(n768), .B2(n3177), .ZN(n1381) );
  OAI22_X1 U659 ( .A1(n3173), .A2(n2243), .B1(n765), .B2(n3177), .ZN(n1378) );
  OAI22_X1 U660 ( .A1(n3173), .A2(n2235), .B1(n771), .B2(n3176), .ZN(n1384) );
  OAI22_X1 U661 ( .A1(n3173), .A2(n2245), .B1(n764), .B2(n3177), .ZN(n1377) );
  OAI22_X1 U662 ( .A1(n3173), .A2(n2233), .B1(n772), .B2(n3176), .ZN(n1385) );
  OAI22_X1 U663 ( .A1(n3173), .A2(n2248), .B1(n763), .B2(n3178), .ZN(n1376) );
  OAI22_X1 U664 ( .A1(n3173), .A2(n2231), .B1(n773), .B2(n3176), .ZN(n1386) );
  OAI22_X1 U665 ( .A1(n3173), .A2(n2250), .B1(n762), .B2(n3178), .ZN(n1375) );
  OAI22_X1 U666 ( .A1(n3173), .A2(n2229), .B1(n774), .B2(n3176), .ZN(n1387) );
  OAI22_X1 U667 ( .A1(n3173), .A2(n2252), .B1(n761), .B2(n3178), .ZN(n1374) );
  OAI22_X1 U668 ( .A1(n3172), .A2(n2227), .B1(n775), .B2(n3175), .ZN(n1388) );
  OAI22_X1 U669 ( .A1(n3173), .A2(n2254), .B1(n760), .B2(n3178), .ZN(n1373) );
  OAI22_X1 U670 ( .A1(n3173), .A2(n2225), .B1(n776), .B2(n3175), .ZN(n1389) );
  OAI22_X1 U671 ( .A1(n3172), .A2(n2223), .B1(n777), .B2(n3175), .ZN(n1390) );
  OAI22_X1 U672 ( .A1(n3172), .A2(n2221), .B1(n778), .B2(n3177), .ZN(n1391) );
  OAI22_X1 U673 ( .A1(n3173), .A2(n2260), .B1(n757), .B2(n3179), .ZN(n1370) );
  OAI22_X1 U674 ( .A1(n3172), .A2(n2219), .B1(n779), .B2(n3175), .ZN(n1392) );
  OAI22_X1 U675 ( .A1(n3172), .A2(n2217), .B1(n780), .B2(n3174), .ZN(n1393) );
  OAI22_X1 U676 ( .A1(n3172), .A2(n2215), .B1(n781), .B2(n3174), .ZN(n1394) );
  OAI22_X1 U677 ( .A1(n3173), .A2(n2266), .B1(n754), .B2(n3180), .ZN(n1367) );
  OAI22_X1 U678 ( .A1(n3172), .A2(n2213), .B1(n782), .B2(n3174), .ZN(n1395) );
  OAI22_X1 U679 ( .A1(n3172), .A2(n2268), .B1(n753), .B2(n3180), .ZN(n1366) );
  OAI22_X1 U680 ( .A1(n3172), .A2(n2210), .B1(n783), .B2(n3174), .ZN(n1396) );
  OAI22_X1 U681 ( .A1(n3173), .A2(n2256), .B1(n759), .B2(n3179), .ZN(n1372) );
  OAI22_X1 U682 ( .A1(n3173), .A2(n2258), .B1(n758), .B2(n3179), .ZN(n1371) );
  OAI22_X1 U683 ( .A1(n3173), .A2(n2262), .B1(n756), .B2(n3179), .ZN(n1369) );
  OAI22_X1 U684 ( .A1(n3173), .A2(n2264), .B1(n755), .B2(n3180), .ZN(n1368) );
  OAI22_X1 U685 ( .A1(n2235), .A2(n2973), .B1(n803), .B2(n3110), .ZN(n1416) );
  OAI22_X1 U686 ( .A1(n2250), .A2(n2973), .B1(n793), .B2(n3110), .ZN(n1406) );
  OAI22_X1 U687 ( .A1(n2256), .A2(n2974), .B1(n790), .B2(n3110), .ZN(n1403) );
  OAI22_X1 U688 ( .A1(n2221), .A2(n2972), .B1(n810), .B2(n3110), .ZN(n1423) );
  OAI22_X1 U689 ( .A1(n2262), .A2(n2974), .B1(n787), .B2(n3110), .ZN(n1400) );
  OAI22_X1 U690 ( .A1(n2235), .A2(n2979), .B1(n867), .B2(n3120), .ZN(n1480) );
  OAI22_X1 U691 ( .A1(n2250), .A2(n2979), .B1(n857), .B2(n3120), .ZN(n1470) );
  OAI22_X1 U692 ( .A1(n2256), .A2(n2980), .B1(n854), .B2(n3120), .ZN(n1467) );
  OAI22_X1 U693 ( .A1(n2221), .A2(n2978), .B1(n874), .B2(n3120), .ZN(n1487) );
  OAI22_X1 U694 ( .A1(n2262), .A2(n2980), .B1(n851), .B2(n3120), .ZN(n1464) );
  OAI22_X1 U695 ( .A1(n2213), .A2(n2975), .B1(n846), .B2(n3115), .ZN(n1459) );
  OAI22_X1 U696 ( .A1(n2243), .A2(n2976), .B1(n828), .B2(n3115), .ZN(n1441) );
  OAI22_X1 U697 ( .A1(n2235), .A2(n2985), .B1(n931), .B2(n3130), .ZN(n1544) );
  OAI22_X1 U698 ( .A1(n2250), .A2(n2985), .B1(n921), .B2(n3130), .ZN(n1534) );
  OAI22_X1 U699 ( .A1(n2256), .A2(n2986), .B1(n918), .B2(n3130), .ZN(n1531) );
  OAI22_X1 U700 ( .A1(n2221), .A2(n2984), .B1(n938), .B2(n3130), .ZN(n1551) );
  OAI22_X1 U701 ( .A1(n2260), .A2(n2977), .B1(n820), .B2(n3115), .ZN(n1433) );
  OAI22_X1 U702 ( .A1(n2262), .A2(n2977), .B1(n819), .B2(n3115), .ZN(n1432) );
  OAI22_X1 U703 ( .A1(n2262), .A2(n2986), .B1(n915), .B2(n3130), .ZN(n1528) );
  OAI22_X1 U704 ( .A1(n2235), .A2(n2982), .B1(n899), .B2(n3125), .ZN(n1512) );
  OAI22_X1 U705 ( .A1(n2221), .A2(n2981), .B1(n906), .B2(n3125), .ZN(n1519) );
  OAI22_X1 U706 ( .A1(n2250), .A2(n2982), .B1(n889), .B2(n3125), .ZN(n1502) );
  OAI22_X1 U707 ( .A1(n2256), .A2(n2983), .B1(n886), .B2(n3125), .ZN(n1499) );
  OAI22_X1 U708 ( .A1(n2262), .A2(n2983), .B1(n883), .B2(n3125), .ZN(n1496) );
  NAND2_X1 U709 ( .A1(n994), .A2(n2335), .ZN(n1607) );
  NAND2_X1 U710 ( .A1(n801), .A2(n2972), .ZN(n1414) );
  NAND2_X1 U711 ( .A1(n797), .A2(n2972), .ZN(n1410) );
  NAND2_X1 U712 ( .A1(n802), .A2(n2972), .ZN(n1415) );
  NAND2_X1 U713 ( .A1(n894), .A2(n2981), .ZN(n1507) );
  NAND2_X1 U714 ( .A1(n897), .A2(n2981), .ZN(n1510) );
  NAND2_X1 U715 ( .A1(n898), .A2(n2981), .ZN(n1511) );
  NAND2_X1 U716 ( .A1(n830), .A2(n2975), .ZN(n1443) );
  NAND2_X1 U717 ( .A1(n829), .A2(n2975), .ZN(n1442) );
  NAND2_X1 U718 ( .A1(n834), .A2(n2975), .ZN(n1447) );
  NAND2_X1 U719 ( .A1(n861), .A2(n2978), .ZN(n1474) );
  NAND2_X1 U720 ( .A1(n866), .A2(n2978), .ZN(n1479) );
  NAND2_X1 U721 ( .A1(n929), .A2(n2984), .ZN(n1542) );
  NAND2_X1 U722 ( .A1(n930), .A2(n2984), .ZN(n1543) );
  NAND2_X1 U723 ( .A1(n958), .A2(n2987), .ZN(n1571) );
  NAND2_X1 U724 ( .A1(n962), .A2(n2987), .ZN(n1575) );
  INV_X1 U725 ( .A(n2484), .ZN(PRED[1]) );
  AOI222_X1 U726 ( .A1(PRED_TK[1]), .A2(n2462), .B1(NEXT_PC[1]), .B2(n3093), 
        .C1(NEW_PC[1]), .C2(n3102), .ZN(n2484) );
  INV_X1 U727 ( .A(n2066), .ZN(n1861) );
  AOI22_X1 U728 ( .A1(n3168), .A2(n373), .B1(n2053), .B2(CURR_PC[1]), .ZN(
        n2066) );
  INV_X1 U729 ( .A(n2068), .ZN(n1857) );
  AOI22_X1 U730 ( .A1(n3168), .A2(n453), .B1(n2053), .B2(CURR_PC[6]), .ZN(
        n2068) );
  INV_X1 U731 ( .A(n2065), .ZN(n1864) );
  AOI22_X1 U732 ( .A1(n3167), .A2(n469), .B1(n2053), .B2(CURR_PC[7]), .ZN(
        n2065) );
  INV_X1 U733 ( .A(n2069), .ZN(n1856) );
  AOI22_X1 U734 ( .A1(n3168), .A2(n485), .B1(n2053), .B2(CURR_PC[8]), .ZN(
        n2069) );
  INV_X1 U735 ( .A(n2064), .ZN(n1865) );
  AOI22_X1 U736 ( .A1(n3168), .A2(n501), .B1(n2053), .B2(CURR_PC[9]), .ZN(
        n2064) );
  INV_X1 U737 ( .A(n2070), .ZN(n1855) );
  AOI22_X1 U738 ( .A1(n3167), .A2(n517), .B1(n2053), .B2(CURR_PC[10]), .ZN(
        n2070) );
  INV_X1 U739 ( .A(n2063), .ZN(n1866) );
  AOI22_X1 U740 ( .A1(n3168), .A2(n533), .B1(n2053), .B2(CURR_PC[11]), .ZN(
        n2063) );
  INV_X1 U741 ( .A(n2071), .ZN(n1854) );
  AOI22_X1 U742 ( .A1(n3167), .A2(n549), .B1(n2053), .B2(CURR_PC[12]), .ZN(
        n2071) );
  INV_X1 U743 ( .A(n2062), .ZN(n1867) );
  AOI22_X1 U744 ( .A1(n3167), .A2(n565), .B1(n2053), .B2(CURR_PC[13]), .ZN(
        n2062) );
  INV_X1 U745 ( .A(n2060), .ZN(n1869) );
  AOI22_X1 U746 ( .A1(n3167), .A2(n629), .B1(n2053), .B2(CURR_PC[17]), .ZN(
        n2060) );
  INV_X1 U747 ( .A(n2051), .ZN(n1876) );
  AOI22_X1 U748 ( .A1(n3167), .A2(n341), .B1(n2053), .B2(CURR_PC[31]), .ZN(
        n2051) );
  INV_X1 U749 ( .A(n2072), .ZN(n1853) );
  AOI22_X1 U750 ( .A1(n3167), .A2(n581), .B1(n2053), .B2(CURR_PC[14]), .ZN(
        n2072) );
  INV_X1 U751 ( .A(n2061), .ZN(n1868) );
  AOI22_X1 U752 ( .A1(n2052), .A2(n597), .B1(n2053), .B2(CURR_PC[15]), .ZN(
        n2061) );
  INV_X1 U753 ( .A(n2073), .ZN(n1852) );
  AOI22_X1 U754 ( .A1(n3167), .A2(n613), .B1(n2053), .B2(CURR_PC[16]), .ZN(
        n2073) );
  INV_X1 U755 ( .A(n2074), .ZN(n1851) );
  AOI22_X1 U756 ( .A1(n2052), .A2(n645), .B1(n2053), .B2(CURR_PC[18]), .ZN(
        n2074) );
  INV_X1 U757 ( .A(n2059), .ZN(n1870) );
  AOI22_X1 U758 ( .A1(n3168), .A2(n661), .B1(n2053), .B2(CURR_PC[19]), .ZN(
        n2059) );
  INV_X1 U759 ( .A(n2075), .ZN(n1850) );
  AOI22_X1 U760 ( .A1(n2052), .A2(n677), .B1(n2053), .B2(CURR_PC[20]), .ZN(
        n2075) );
  INV_X1 U761 ( .A(n2058), .ZN(n1871) );
  AOI22_X1 U762 ( .A1(n2052), .A2(n699), .B1(n2053), .B2(CURR_PC[21]), .ZN(
        n2058) );
  INV_X1 U763 ( .A(n2076), .ZN(n1849) );
  AOI22_X1 U764 ( .A1(n3167), .A2(n197), .B1(n2053), .B2(CURR_PC[22]), .ZN(
        n2076) );
  INV_X1 U765 ( .A(n2057), .ZN(n1872) );
  AOI22_X1 U766 ( .A1(n2052), .A2(n213), .B1(n2053), .B2(CURR_PC[23]), .ZN(
        n2057) );
  INV_X1 U767 ( .A(n2077), .ZN(n1848) );
  AOI22_X1 U768 ( .A1(n3168), .A2(n229), .B1(n2053), .B2(CURR_PC[24]), .ZN(
        n2077) );
  INV_X1 U769 ( .A(n2056), .ZN(n1873) );
  AOI22_X1 U770 ( .A1(n2052), .A2(n245), .B1(n2053), .B2(CURR_PC[25]), .ZN(
        n2056) );
  INV_X1 U771 ( .A(n2078), .ZN(n1847) );
  AOI22_X1 U772 ( .A1(n3168), .A2(n261), .B1(n2053), .B2(CURR_PC[26]), .ZN(
        n2078) );
  INV_X1 U773 ( .A(n2055), .ZN(n1874) );
  AOI22_X1 U774 ( .A1(n2052), .A2(n277), .B1(n2053), .B2(CURR_PC[27]), .ZN(
        n2055) );
  INV_X1 U775 ( .A(n2079), .ZN(n1846) );
  AOI22_X1 U776 ( .A1(n2052), .A2(n293), .B1(n2053), .B2(CURR_PC[28]), .ZN(
        n2079) );
  INV_X1 U777 ( .A(n2054), .ZN(n1875) );
  AOI22_X1 U778 ( .A1(n3168), .A2(n309), .B1(n2053), .B2(CURR_PC[29]), .ZN(
        n2054) );
  INV_X1 U779 ( .A(n2080), .ZN(n1845) );
  AOI22_X1 U780 ( .A1(n3167), .A2(n325), .B1(n2053), .B2(CURR_PC[30]), .ZN(
        n2080) );
  INV_X1 U781 ( .A(n2164), .ZN(n1760) );
  AOI22_X1 U782 ( .A1(CURR_PC[8]), .A2(n3159), .B1(n2148), .B2(n1411), .ZN(
        n2164) );
  INV_X1 U783 ( .A(n2159), .ZN(n1769) );
  AOI22_X1 U784 ( .A1(CURR_PC[9]), .A2(n3159), .B1(n2148), .B2(n1446), .ZN(
        n2159) );
  INV_X1 U785 ( .A(n2165), .ZN(n1759) );
  AOI22_X1 U786 ( .A1(CURR_PC[10]), .A2(n3157), .B1(n2148), .B2(n1475), .ZN(
        n2165) );
  INV_X1 U787 ( .A(n2167), .ZN(n1757) );
  AOI22_X1 U788 ( .A1(CURR_PC[14]), .A2(n3157), .B1(n2148), .B2(n1478), .ZN(
        n2167) );
  INV_X1 U789 ( .A(n2151), .ZN(n1777) );
  AOI22_X1 U790 ( .A1(CURR_PC[25]), .A2(n3157), .B1(n2148), .B2(n1506), .ZN(
        n2151) );
  INV_X1 U791 ( .A(n2149), .ZN(n1779) );
  AOI22_X1 U792 ( .A1(CURR_PC[29]), .A2(n3157), .B1(n2148), .B2(n1538), .ZN(
        n2149) );
  INV_X1 U793 ( .A(n2175), .ZN(n1749) );
  AOI22_X1 U794 ( .A1(CURR_PC[30]), .A2(n3159), .B1(n2148), .B2(n1539), .ZN(
        n2175) );
  INV_X1 U795 ( .A(n2146), .ZN(n1780) );
  AOI22_X1 U796 ( .A1(CURR_PC[31]), .A2(n3159), .B1(n2148), .B2(n1570), .ZN(
        n2146) );
  INV_X1 U797 ( .A(n2161), .ZN(n1765) );
  AOI22_X1 U798 ( .A1(CURR_PC[1]), .A2(n3159), .B1(n2148), .B2(n1795), .ZN(
        n2161) );
  INV_X1 U799 ( .A(n2160), .ZN(n1768) );
  AOI22_X1 U800 ( .A1(CURR_PC[7]), .A2(n3160), .B1(n2148), .B2(n1799), .ZN(
        n2160) );
  INV_X1 U801 ( .A(n2158), .ZN(n1770) );
  AOI22_X1 U802 ( .A1(CURR_PC[11]), .A2(n3160), .B1(n2148), .B2(n1826), .ZN(
        n2158) );
  INV_X1 U803 ( .A(n2166), .ZN(n1758) );
  AOI22_X1 U804 ( .A1(CURR_PC[12]), .A2(n3160), .B1(n2148), .B2(n1830), .ZN(
        n2166) );
  INV_X1 U805 ( .A(n2150), .ZN(n1778) );
  AOI22_X1 U806 ( .A1(CURR_PC[27]), .A2(n3160), .B1(n2148), .B2(n1831), .ZN(
        n2150) );
  INV_X1 U807 ( .A(n2174), .ZN(n1750) );
  AOI22_X1 U808 ( .A1(CURR_PC[28]), .A2(n3160), .B1(n2148), .B2(n1858), .ZN(
        n2174) );
  INV_X1 U809 ( .A(n2162), .ZN(n1764) );
  AOI22_X1 U810 ( .A1(CURR_PC[0]), .A2(n3158), .B1(n2148), .B2(n1885), .ZN(
        n2162) );
  INV_X1 U811 ( .A(n2163), .ZN(n1761) );
  AOI22_X1 U812 ( .A1(CURR_PC[6]), .A2(n3158), .B1(n2148), .B2(n1886), .ZN(
        n2163) );
  INV_X1 U813 ( .A(n2157), .ZN(n1771) );
  AOI22_X1 U814 ( .A1(CURR_PC[13]), .A2(n3157), .B1(n2148), .B2(n1887), .ZN(
        n2157) );
  INV_X1 U815 ( .A(n2156), .ZN(n1772) );
  AOI22_X1 U816 ( .A1(CURR_PC[15]), .A2(n3157), .B1(n2148), .B2(n1888), .ZN(
        n2156) );
  INV_X1 U817 ( .A(n2168), .ZN(n1756) );
  AOI22_X1 U818 ( .A1(CURR_PC[16]), .A2(n3158), .B1(n2148), .B2(n1889), .ZN(
        n2168) );
  INV_X1 U819 ( .A(n2155), .ZN(n1773) );
  AOI22_X1 U820 ( .A1(CURR_PC[17]), .A2(n3160), .B1(n2148), .B2(n1890), .ZN(
        n2155) );
  INV_X1 U821 ( .A(n2169), .ZN(n1755) );
  AOI22_X1 U822 ( .A1(CURR_PC[18]), .A2(n3159), .B1(n2148), .B2(n1891), .ZN(
        n2169) );
  INV_X1 U823 ( .A(n2154), .ZN(n1774) );
  AOI22_X1 U824 ( .A1(CURR_PC[19]), .A2(n3158), .B1(n2148), .B2(n1892), .ZN(
        n2154) );
  INV_X1 U825 ( .A(n2153), .ZN(n1775) );
  AOI22_X1 U826 ( .A1(CURR_PC[21]), .A2(n3159), .B1(n2148), .B2(n1893), .ZN(
        n2153) );
  INV_X1 U827 ( .A(n2152), .ZN(n1776) );
  AOI22_X1 U828 ( .A1(CURR_PC[23]), .A2(n3158), .B1(n2148), .B2(n1894), .ZN(
        n2152) );
  INV_X1 U829 ( .A(n2170), .ZN(n1754) );
  AOI22_X1 U830 ( .A1(CURR_PC[20]), .A2(n3158), .B1(n2148), .B2(n1940), .ZN(
        n2170) );
  INV_X1 U831 ( .A(n2171), .ZN(n1753) );
  AOI22_X1 U832 ( .A1(CURR_PC[22]), .A2(n3160), .B1(n2148), .B2(n1941), .ZN(
        n2171) );
  INV_X1 U833 ( .A(n2172), .ZN(n1752) );
  AOI22_X1 U834 ( .A1(CURR_PC[24]), .A2(n3157), .B1(n2148), .B2(n1942), .ZN(
        n2172) );
  INV_X1 U835 ( .A(n2173), .ZN(n1751) );
  AOI22_X1 U836 ( .A1(CURR_PC[26]), .A2(n3157), .B1(n2148), .B2(n1943), .ZN(
        n2173) );
  INV_X1 U837 ( .A(n2098), .ZN(n1829) );
  AOI22_X1 U838 ( .A1(n2084), .A2(n374), .B1(CURR_PC[1]), .B2(n3165), .ZN(
        n2098) );
  INV_X1 U839 ( .A(n2100), .ZN(n1825) );
  AOI22_X1 U840 ( .A1(n2084), .A2(n454), .B1(CURR_PC[6]), .B2(n3164), .ZN(
        n2100) );
  INV_X1 U841 ( .A(n2097), .ZN(n1832) );
  AOI22_X1 U842 ( .A1(n2084), .A2(n470), .B1(CURR_PC[7]), .B2(n3166), .ZN(
        n2097) );
  INV_X1 U843 ( .A(n2101), .ZN(n1824) );
  AOI22_X1 U844 ( .A1(n2084), .A2(n486), .B1(CURR_PC[8]), .B2(n3165), .ZN(
        n2101) );
  INV_X1 U845 ( .A(n2096), .ZN(n1833) );
  AOI22_X1 U846 ( .A1(n2084), .A2(n502), .B1(CURR_PC[9]), .B2(n3166), .ZN(
        n2096) );
  INV_X1 U847 ( .A(n2102), .ZN(n1823) );
  AOI22_X1 U848 ( .A1(n2084), .A2(n518), .B1(CURR_PC[10]), .B2(n3164), .ZN(
        n2102) );
  INV_X1 U849 ( .A(n2103), .ZN(n1822) );
  AOI22_X1 U850 ( .A1(n2084), .A2(n550), .B1(CURR_PC[12]), .B2(n3163), .ZN(
        n2103) );
  INV_X1 U851 ( .A(n2094), .ZN(n1835) );
  AOI22_X1 U852 ( .A1(n2084), .A2(n566), .B1(CURR_PC[13]), .B2(n3166), .ZN(
        n2094) );
  INV_X1 U853 ( .A(n2104), .ZN(n1821) );
  AOI22_X1 U854 ( .A1(n2084), .A2(n582), .B1(CURR_PC[14]), .B2(n3166), .ZN(
        n2104) );
  INV_X1 U855 ( .A(n2088), .ZN(n1841) );
  AOI22_X1 U856 ( .A1(n2084), .A2(n246), .B1(CURR_PC[25]), .B2(n3166), .ZN(
        n2088) );
  INV_X1 U857 ( .A(n2083), .ZN(n1844) );
  AOI22_X1 U858 ( .A1(n2084), .A2(n342), .B1(CURR_PC[31]), .B2(n3165), .ZN(
        n2083) );
  INV_X1 U859 ( .A(n2099), .ZN(n1828) );
  AOI22_X1 U860 ( .A1(n2084), .A2(n358), .B1(CURR_PC[0]), .B2(n3165), .ZN(
        n2099) );
  INV_X1 U861 ( .A(n2095), .ZN(n1834) );
  AOI22_X1 U862 ( .A1(n2084), .A2(n534), .B1(CURR_PC[11]), .B2(n3163), .ZN(
        n2095) );
  INV_X1 U863 ( .A(n2093), .ZN(n1836) );
  AOI22_X1 U864 ( .A1(n2084), .A2(n598), .B1(CURR_PC[15]), .B2(n3163), .ZN(
        n2093) );
  INV_X1 U865 ( .A(n2092), .ZN(n1837) );
  AOI22_X1 U866 ( .A1(n2084), .A2(n630), .B1(CURR_PC[17]), .B2(n3164), .ZN(
        n2092) );
  INV_X1 U867 ( .A(n2091), .ZN(n1838) );
  AOI22_X1 U868 ( .A1(n2084), .A2(n662), .B1(CURR_PC[19]), .B2(n3165), .ZN(
        n2091) );
  INV_X1 U869 ( .A(n2090), .ZN(n1839) );
  AOI22_X1 U870 ( .A1(n2084), .A2(n700), .B1(CURR_PC[21]), .B2(n3163), .ZN(
        n2090) );
  INV_X1 U871 ( .A(n2089), .ZN(n1840) );
  AOI22_X1 U872 ( .A1(n2084), .A2(n214), .B1(CURR_PC[23]), .B2(n3164), .ZN(
        n2089) );
  INV_X1 U873 ( .A(n2087), .ZN(n1842) );
  AOI22_X1 U874 ( .A1(n2084), .A2(n278), .B1(CURR_PC[27]), .B2(n3163), .ZN(
        n2087) );
  INV_X1 U875 ( .A(n2086), .ZN(n1843) );
  AOI22_X1 U876 ( .A1(n2084), .A2(n310), .B1(CURR_PC[29]), .B2(n3164), .ZN(
        n2086) );
  INV_X1 U877 ( .A(n2112), .ZN(n1813) );
  AOI22_X1 U878 ( .A1(n2084), .A2(n326), .B1(CURR_PC[30]), .B2(n3166), .ZN(
        n2112) );
  INV_X1 U879 ( .A(n2105), .ZN(n1820) );
  AOI22_X1 U880 ( .A1(n2084), .A2(n614), .B1(CURR_PC[16]), .B2(n3164), .ZN(
        n2105) );
  INV_X1 U881 ( .A(n2106), .ZN(n1819) );
  AOI22_X1 U882 ( .A1(n2084), .A2(n646), .B1(CURR_PC[18]), .B2(n3163), .ZN(
        n2106) );
  INV_X1 U883 ( .A(n2107), .ZN(n1818) );
  AOI22_X1 U884 ( .A1(n2084), .A2(n678), .B1(CURR_PC[20]), .B2(n3165), .ZN(
        n2107) );
  INV_X1 U885 ( .A(n2108), .ZN(n1817) );
  AOI22_X1 U886 ( .A1(n2084), .A2(n198), .B1(CURR_PC[22]), .B2(n3164), .ZN(
        n2108) );
  INV_X1 U887 ( .A(n2109), .ZN(n1816) );
  AOI22_X1 U888 ( .A1(n2084), .A2(n230), .B1(CURR_PC[24]), .B2(n3163), .ZN(
        n2109) );
  INV_X1 U889 ( .A(n2110), .ZN(n1815) );
  AOI22_X1 U890 ( .A1(n2084), .A2(n262), .B1(CURR_PC[26]), .B2(n3166), .ZN(
        n2110) );
  INV_X1 U891 ( .A(n2111), .ZN(n1814) );
  AOI22_X1 U892 ( .A1(n2084), .A2(n294), .B1(CURR_PC[28]), .B2(n3163), .ZN(
        n2111) );
  OR2_X1 U893 ( .A1(n1918), .A2(n2116), .ZN(n1798) );
  OR2_X1 U894 ( .A1(n418), .A2(n2179), .ZN(n1730) );
  INV_X1 U895 ( .A(n2067), .ZN(n1860) );
  AOI22_X1 U896 ( .A1(n3168), .A2(n357), .B1(CURR_PC[0]), .B2(n2053), .ZN(
        n2067) );
  INV_X1 U897 ( .A(n2193), .ZN(n1732) );
  AOI22_X1 U898 ( .A1(n3155), .A2(n354), .B1(CURR_PC[0]), .B2(n2179), .ZN(
        n2193) );
  INV_X1 U899 ( .A(n2192), .ZN(n1733) );
  AOI22_X1 U900 ( .A1(n3156), .A2(n370), .B1(CURR_PC[1]), .B2(n2179), .ZN(
        n2192) );
  INV_X1 U901 ( .A(n2131), .ZN(n1796) );
  AOI22_X1 U902 ( .A1(CURR_PC[0]), .A2(n2116), .B1(n3162), .B2(n137), .ZN(
        n2131) );
  INV_X1 U903 ( .A(n2130), .ZN(n1797) );
  AOI22_X1 U904 ( .A1(CURR_PC[1]), .A2(n2116), .B1(n3162), .B2(n138), .ZN(
        n2130) );
  INV_X1 U905 ( .A(n2194), .ZN(n1729) );
  AOI22_X1 U906 ( .A1(n3156), .A2(n450), .B1(CURR_PC[6]), .B2(n2179), .ZN(
        n2194) );
  INV_X1 U907 ( .A(n2191), .ZN(n1736) );
  AOI22_X1 U908 ( .A1(n3155), .A2(n466), .B1(CURR_PC[7]), .B2(n2179), .ZN(
        n2191) );
  INV_X1 U909 ( .A(n2195), .ZN(n1728) );
  AOI22_X1 U910 ( .A1(n3156), .A2(n482), .B1(CURR_PC[8]), .B2(n2179), .ZN(
        n2195) );
  INV_X1 U911 ( .A(n2190), .ZN(n1737) );
  AOI22_X1 U912 ( .A1(n3155), .A2(n498), .B1(CURR_PC[9]), .B2(n2179), .ZN(
        n2190) );
  INV_X1 U913 ( .A(n2196), .ZN(n1727) );
  AOI22_X1 U914 ( .A1(n3156), .A2(n514), .B1(CURR_PC[10]), .B2(n2179), .ZN(
        n2196) );
  INV_X1 U915 ( .A(n2197), .ZN(n1726) );
  AOI22_X1 U916 ( .A1(n2178), .A2(n546), .B1(CURR_PC[12]), .B2(n2179), .ZN(
        n2197) );
  INV_X1 U917 ( .A(n2188), .ZN(n1739) );
  AOI22_X1 U918 ( .A1(n3156), .A2(n562), .B1(CURR_PC[13]), .B2(n2179), .ZN(
        n2188) );
  INV_X1 U919 ( .A(n2198), .ZN(n1725) );
  AOI22_X1 U920 ( .A1(n3155), .A2(n578), .B1(CURR_PC[14]), .B2(n2179), .ZN(
        n2198) );
  INV_X1 U921 ( .A(n2182), .ZN(n1745) );
  AOI22_X1 U922 ( .A1(n2178), .A2(n242), .B1(CURR_PC[25]), .B2(n2179), .ZN(
        n2182) );
  INV_X1 U923 ( .A(n2177), .ZN(n1748) );
  AOI22_X1 U924 ( .A1(n3156), .A2(n338), .B1(CURR_PC[31]), .B2(n2179), .ZN(
        n2177) );
  INV_X1 U925 ( .A(n2189), .ZN(n1738) );
  AOI22_X1 U926 ( .A1(n3155), .A2(n530), .B1(CURR_PC[11]), .B2(n2179), .ZN(
        n2189) );
  INV_X1 U927 ( .A(n2187), .ZN(n1740) );
  AOI22_X1 U928 ( .A1(n3155), .A2(n594), .B1(CURR_PC[15]), .B2(n2179), .ZN(
        n2187) );
  INV_X1 U929 ( .A(n2186), .ZN(n1741) );
  AOI22_X1 U930 ( .A1(n3155), .A2(n626), .B1(CURR_PC[17]), .B2(n2179), .ZN(
        n2186) );
  INV_X1 U931 ( .A(n2185), .ZN(n1742) );
  AOI22_X1 U932 ( .A1(n2178), .A2(n658), .B1(CURR_PC[19]), .B2(n2179), .ZN(
        n2185) );
  INV_X1 U933 ( .A(n2184), .ZN(n1743) );
  AOI22_X1 U934 ( .A1(n3155), .A2(n690), .B1(CURR_PC[21]), .B2(n2179), .ZN(
        n2184) );
  INV_X1 U935 ( .A(n2183), .ZN(n1744) );
  AOI22_X1 U936 ( .A1(n3156), .A2(n210), .B1(CURR_PC[23]), .B2(n2179), .ZN(
        n2183) );
  INV_X1 U937 ( .A(n2181), .ZN(n1746) );
  AOI22_X1 U938 ( .A1(n2178), .A2(n274), .B1(CURR_PC[27]), .B2(n2179), .ZN(
        n2181) );
  INV_X1 U939 ( .A(n2180), .ZN(n1747) );
  AOI22_X1 U940 ( .A1(n3156), .A2(n306), .B1(CURR_PC[29]), .B2(n2179), .ZN(
        n2180) );
  INV_X1 U941 ( .A(n2206), .ZN(n1717) );
  AOI22_X1 U942 ( .A1(n2178), .A2(n322), .B1(CURR_PC[30]), .B2(n2179), .ZN(
        n2206) );
  INV_X1 U943 ( .A(n2199), .ZN(n1724) );
  AOI22_X1 U944 ( .A1(n2178), .A2(n610), .B1(CURR_PC[16]), .B2(n2179), .ZN(
        n2199) );
  INV_X1 U945 ( .A(n2200), .ZN(n1723) );
  AOI22_X1 U946 ( .A1(n3156), .A2(n642), .B1(CURR_PC[18]), .B2(n2179), .ZN(
        n2200) );
  INV_X1 U947 ( .A(n2201), .ZN(n1722) );
  AOI22_X1 U948 ( .A1(n3155), .A2(n674), .B1(CURR_PC[20]), .B2(n2179), .ZN(
        n2201) );
  INV_X1 U949 ( .A(n2202), .ZN(n1721) );
  AOI22_X1 U950 ( .A1(n2178), .A2(n194), .B1(CURR_PC[22]), .B2(n2179), .ZN(
        n2202) );
  INV_X1 U951 ( .A(n2203), .ZN(n1720) );
  AOI22_X1 U952 ( .A1(n2178), .A2(n226), .B1(CURR_PC[24]), .B2(n2179), .ZN(
        n2203) );
  INV_X1 U953 ( .A(n2204), .ZN(n1719) );
  AOI22_X1 U954 ( .A1(n3156), .A2(n258), .B1(CURR_PC[26]), .B2(n2179), .ZN(
        n2204) );
  INV_X1 U955 ( .A(n2205), .ZN(n1718) );
  AOI22_X1 U956 ( .A1(n3155), .A2(n290), .B1(CURR_PC[28]), .B2(n2179), .ZN(
        n2205) );
  INV_X1 U957 ( .A(n2132), .ZN(n1793) );
  AOI22_X1 U958 ( .A1(CURR_PC[6]), .A2(n2116), .B1(n3162), .B2(n3), .ZN(n2132)
         );
  INV_X1 U959 ( .A(n2133), .ZN(n1792) );
  AOI22_X1 U960 ( .A1(CURR_PC[8]), .A2(n2116), .B1(n3162), .B2(n4), .ZN(n2133)
         );
  INV_X1 U961 ( .A(n2134), .ZN(n1791) );
  AOI22_X1 U962 ( .A1(CURR_PC[10]), .A2(n2116), .B1(n3161), .B2(n5), .ZN(n2134) );
  INV_X1 U963 ( .A(n2125), .ZN(n1804) );
  AOI22_X1 U964 ( .A1(CURR_PC[15]), .A2(n2116), .B1(n3161), .B2(n6), .ZN(n2125) );
  INV_X1 U965 ( .A(n2124), .ZN(n1805) );
  AOI22_X1 U966 ( .A1(CURR_PC[17]), .A2(n2116), .B1(n3161), .B2(n7), .ZN(n2124) );
  INV_X1 U967 ( .A(n2123), .ZN(n1806) );
  AOI22_X1 U968 ( .A1(CURR_PC[19]), .A2(n2116), .B1(n3161), .B2(n9), .ZN(n2123) );
  INV_X1 U969 ( .A(n2141), .ZN(n1784) );
  AOI22_X1 U970 ( .A1(CURR_PC[24]), .A2(n2116), .B1(n2117), .B2(n42), .ZN(
        n2141) );
  INV_X1 U971 ( .A(n2142), .ZN(n1783) );
  AOI22_X1 U972 ( .A1(CURR_PC[26]), .A2(n2116), .B1(n3161), .B2(n43), .ZN(
        n2142) );
  INV_X1 U973 ( .A(n2143), .ZN(n1782) );
  AOI22_X1 U974 ( .A1(CURR_PC[28]), .A2(n2116), .B1(n3161), .B2(n44), .ZN(
        n2143) );
  INV_X1 U975 ( .A(n2128), .ZN(n1801) );
  AOI22_X1 U976 ( .A1(CURR_PC[9]), .A2(n2116), .B1(n2117), .B2(n52), .ZN(n2128) );
  INV_X1 U977 ( .A(n2127), .ZN(n1802) );
  AOI22_X1 U978 ( .A1(CURR_PC[11]), .A2(n2116), .B1(n3162), .B2(n55), .ZN(
        n2127) );
  INV_X1 U979 ( .A(n2135), .ZN(n1790) );
  AOI22_X1 U980 ( .A1(CURR_PC[12]), .A2(n2116), .B1(n3161), .B2(n56), .ZN(
        n2135) );
  INV_X1 U981 ( .A(n2126), .ZN(n1803) );
  AOI22_X1 U982 ( .A1(CURR_PC[13]), .A2(n2116), .B1(n3161), .B2(n58), .ZN(
        n2126) );
  INV_X1 U983 ( .A(n2136), .ZN(n1789) );
  AOI22_X1 U984 ( .A1(CURR_PC[14]), .A2(n2116), .B1(n3162), .B2(n59), .ZN(
        n2136) );
  INV_X1 U985 ( .A(n2137), .ZN(n1788) );
  AOI22_X1 U986 ( .A1(CURR_PC[16]), .A2(n2116), .B1(n3162), .B2(n61), .ZN(
        n2137) );
  INV_X1 U987 ( .A(n2119), .ZN(n1810) );
  AOI22_X1 U988 ( .A1(CURR_PC[27]), .A2(n2116), .B1(n2117), .B2(n88), .ZN(
        n2119) );
  INV_X1 U989 ( .A(n2118), .ZN(n1811) );
  AOI22_X1 U990 ( .A1(CURR_PC[29]), .A2(n2116), .B1(n3162), .B2(n89), .ZN(
        n2118) );
  INV_X1 U991 ( .A(n2144), .ZN(n1781) );
  AOI22_X1 U992 ( .A1(CURR_PC[30]), .A2(n2116), .B1(n2117), .B2(n92), .ZN(
        n2144) );
  INV_X1 U993 ( .A(n2115), .ZN(n1812) );
  AOI22_X1 U994 ( .A1(CURR_PC[31]), .A2(n2116), .B1(n3162), .B2(n96), .ZN(
        n2115) );
  INV_X1 U995 ( .A(n2129), .ZN(n1800) );
  AOI22_X1 U996 ( .A1(CURR_PC[7]), .A2(n2116), .B1(n2117), .B2(n139), .ZN(
        n2129) );
  INV_X1 U997 ( .A(n2138), .ZN(n1787) );
  AOI22_X1 U998 ( .A1(CURR_PC[18]), .A2(n2116), .B1(n3161), .B2(n140), .ZN(
        n2138) );
  INV_X1 U999 ( .A(n2139), .ZN(n1786) );
  AOI22_X1 U1000 ( .A1(CURR_PC[20]), .A2(n2116), .B1(n3161), .B2(n141), .ZN(
        n2139) );
  INV_X1 U1001 ( .A(n2122), .ZN(n1807) );
  AOI22_X1 U1002 ( .A1(CURR_PC[21]), .A2(n2116), .B1(n2117), .B2(n142), .ZN(
        n2122) );
  INV_X1 U1003 ( .A(n2140), .ZN(n1785) );
  AOI22_X1 U1004 ( .A1(CURR_PC[22]), .A2(n2116), .B1(n2117), .B2(n143), .ZN(
        n2140) );
  INV_X1 U1005 ( .A(n2121), .ZN(n1808) );
  AOI22_X1 U1006 ( .A1(CURR_PC[23]), .A2(n2116), .B1(n3162), .B2(n144), .ZN(
        n2121) );
  INV_X1 U1007 ( .A(n2120), .ZN(n1809) );
  AOI22_X1 U1008 ( .A1(CURR_PC[25]), .A2(n2116), .B1(n2117), .B2(n145), .ZN(
        n2120) );
  NAND2_X1 U1009 ( .A1(n767), .A2(n3172), .ZN(n1380) );
  NAND2_X1 U1010 ( .A1(n766), .A2(n3172), .ZN(n1379) );
  NAND2_X1 U1011 ( .A1(n769), .A2(n3172), .ZN(n1382) );
  NAND2_X1 U1012 ( .A1(n770), .A2(n3172), .ZN(n1383) );
  INV_X1 U1013 ( .A(n2048), .ZN(n1877) );
  AOI22_X1 U1014 ( .A1(n3180), .A2(CURR_PC[0]), .B1(n3172), .B2(n361), .ZN(
        n2048) );
  OR2_X1 U1015 ( .A1(n1961), .A2(n3159), .ZN(n1766) );
  OR2_X1 U1016 ( .A1(n1960), .A2(n3158), .ZN(n1763) );
  OR2_X1 U1017 ( .A1(n390), .A2(n3164), .ZN(n1827) );
  OR2_X1 U1018 ( .A1(n1958), .A2(n3147), .ZN(n1670) );
  OR2_X1 U1019 ( .A1(n1959), .A2(n3148), .ZN(n1666) );
  NOR2_X1 U1020 ( .A1(n2862), .A2(CURR_PC[3]), .ZN(n2848) );
  NOR2_X1 U1021 ( .A1(CURR_PC[4]), .A2(CURR_PC[5]), .ZN(n2851) );
  AOI221_X1 U1022 ( .B1(n357), .B2(n3085), .C1(n361), .C2(n2504), .A(n2634), 
        .ZN(n2633) );
  OAI22_X1 U1023 ( .A1(n3088), .A2(n2907), .B1(n2332), .B2(n2513), .ZN(n2634)
         );
  AOI221_X1 U1024 ( .B1(n645), .B2(n3086), .C1(n2504), .C2(n2922), .A(n2812), 
        .ZN(n2810) );
  OAI22_X1 U1025 ( .A1(n3087), .A2(n2908), .B1(n3089), .B2(n2514), .ZN(n2812)
         );
  AOI221_X1 U1026 ( .B1(n629), .B2(n2081), .C1(n2504), .C2(n2923), .A(n2801), 
        .ZN(n2799) );
  OAI22_X1 U1027 ( .A1(n3088), .A2(n2909), .B1(n3090), .B2(n2522), .ZN(n2801)
         );
  AOI221_X1 U1028 ( .B1(n597), .B2(n3086), .C1(n2504), .C2(n2924), .A(n2779), 
        .ZN(n2777) );
  OAI22_X1 U1029 ( .A1(n3087), .A2(n2910), .B1(n3089), .B2(n2535), .ZN(n2779)
         );
  AOI221_X1 U1030 ( .B1(n197), .B2(n3086), .C1(n2504), .C2(n2925), .A(n2523), 
        .ZN(n2521) );
  OAI22_X1 U1031 ( .A1(n2269), .A2(n2911), .B1(n3089), .B2(n2546), .ZN(n2523)
         );
  AOI221_X1 U1032 ( .B1(n261), .B2(n3085), .C1(n2504), .C2(n2926), .A(n2569), 
        .ZN(n2567) );
  OAI22_X1 U1033 ( .A1(n3088), .A2(n2912), .B1(n2332), .B2(n2557), .ZN(n2569)
         );
  AOI221_X1 U1034 ( .B1(n325), .B2(n2081), .C1(n2504), .C2(n2927), .A(n2613), 
        .ZN(n2611) );
  OAI22_X1 U1035 ( .A1(n3087), .A2(n2913), .B1(n3090), .B2(n2568), .ZN(n2613)
         );
  AOI221_X1 U1036 ( .B1(n309), .B2(n3085), .C1(n2504), .C2(n2928), .A(n2602), 
        .ZN(n2600) );
  OAI22_X1 U1037 ( .A1(n3088), .A2(n2914), .B1(n2332), .B2(n2579), .ZN(n2602)
         );
  AOI221_X1 U1038 ( .B1(n517), .B2(n3085), .C1(n2504), .C2(n2929), .A(n2724), 
        .ZN(n2722) );
  OAI22_X1 U1039 ( .A1(n2269), .A2(n2915), .B1(n2332), .B2(n2590), .ZN(n2724)
         );
  AOI221_X1 U1040 ( .B1(n581), .B2(n2081), .C1(n2504), .C2(n2930), .A(n2768), 
        .ZN(n2766) );
  OAI22_X1 U1041 ( .A1(n3088), .A2(n2916), .B1(n3090), .B2(n2601), .ZN(n2768)
         );
  AOI221_X1 U1042 ( .B1(n565), .B2(n3085), .C1(n2504), .C2(n2931), .A(n2757), 
        .ZN(n2755) );
  OAI22_X1 U1043 ( .A1(n2269), .A2(n2917), .B1(n2332), .B2(n2612), .ZN(n2757)
         );
  AOI221_X1 U1044 ( .B1(n549), .B2(n3086), .C1(n2504), .C2(n2932), .A(n2746), 
        .ZN(n2744) );
  OAI22_X1 U1045 ( .A1(n3087), .A2(n2918), .B1(n3089), .B2(n2623), .ZN(n2746)
         );
  AOI221_X1 U1046 ( .B1(n341), .B2(n3086), .C1(n2504), .C2(n2952), .A(n2624), 
        .ZN(n2622) );
  OAI22_X1 U1047 ( .A1(n2269), .A2(n2919), .B1(n3089), .B2(n2644), .ZN(n2624)
         );
  AOI221_X1 U1048 ( .B1(n373), .B2(n2081), .C1(n2504), .C2(n2953), .A(n2645), 
        .ZN(n2643) );
  OAI22_X1 U1049 ( .A1(n3087), .A2(n2920), .B1(n3090), .B2(n2653), .ZN(n2645)
         );
  AOI221_X1 U1050 ( .B1(n453), .B2(n3086), .C1(n2504), .C2(n2954), .A(n2680), 
        .ZN(n2678) );
  OAI22_X1 U1051 ( .A1(n3087), .A2(n2921), .B1(n3089), .B2(n2655), .ZN(n2680)
         );
  AOI221_X1 U1052 ( .B1(n2081), .B2(n2950), .C1(n2504), .C2(n2734), .A(n2505), 
        .ZN(n2502) );
  OAI22_X1 U1053 ( .A1(n734), .A2(n3088), .B1(n735), .B2(n2332), .ZN(n2505) );
  OAI22_X1 U1054 ( .A1(n769), .A2(n2372), .B1(n2332), .B2(n2789), .ZN(n2660)
         );
  OAI22_X1 U1055 ( .A1(n1068), .A2(n3081), .B1(n3084), .B2(n2864), .ZN(n2559)
         );
  OAI22_X1 U1056 ( .A1(n1070), .A2(n3080), .B1(n2343), .B2(n2865), .ZN(n2603)
         );
  OAI22_X1 U1057 ( .A1(n3082), .A2(n2866), .B1(n991), .B2(n3083), .ZN(n2635)
         );
  OAI22_X1 U1058 ( .A1(n3080), .A2(n2867), .B1(n983), .B2(n3083), .ZN(n2791)
         );
  OAI22_X1 U1059 ( .A1(n3080), .A2(n2868), .B1(n978), .B2(n3083), .ZN(n2570)
         );
  OAI22_X1 U1060 ( .A1(n3082), .A2(n2869), .B1(n986), .B2(n3083), .ZN(n2725)
         );
  OAI22_X1 U1061 ( .A1(n3082), .A2(n2870), .B1(n995), .B2(n3083), .ZN(n2692)
         );
  OAI22_X1 U1062 ( .A1(n3081), .A2(n2871), .B1(n998), .B2(n3083), .ZN(n2758)
         );
  OAI22_X1 U1063 ( .A1(n743), .A2(n3079), .B1(n742), .B2(n3083), .ZN(n2508) );
  OAI22_X1 U1064 ( .A1(n897), .A2(n3002), .B1(n929), .B2(n2349), .ZN(n2663) );
  OAI22_X1 U1065 ( .A1(n3080), .A2(n2872), .B1(n982), .B2(n2343), .ZN(n2813)
         );
  OAI22_X1 U1066 ( .A1(n3080), .A2(n2873), .B1(n999), .B2(n3084), .ZN(n2780)
         );
  OAI22_X1 U1067 ( .A1(n3082), .A2(n2874), .B1(n980), .B2(n2343), .ZN(n2524)
         );
  OAI22_X1 U1068 ( .A1(n3082), .A2(n2875), .B1(n981), .B2(n3084), .ZN(n2835)
         );
  OAI22_X1 U1069 ( .A1(n3081), .A2(n2876), .B1(n979), .B2(n3084), .ZN(n2548)
         );
  OAI22_X1 U1070 ( .A1(n3080), .A2(n2877), .B1(n976), .B2(n3084), .ZN(n2614)
         );
  OAI22_X1 U1071 ( .A1(n3079), .A2(n2878), .B1(n977), .B2(n2343), .ZN(n2592)
         );
  OAI22_X1 U1072 ( .A1(n3079), .A2(n2879), .B1(n996), .B2(n3084), .ZN(n2714)
         );
  OAI22_X1 U1073 ( .A1(n3080), .A2(n2880), .B1(n987), .B2(n2343), .ZN(n2703)
         );
  OAI22_X1 U1074 ( .A1(n3081), .A2(n2881), .B1(n984), .B2(n2343), .ZN(n2769)
         );
  OAI22_X1 U1075 ( .A1(n3082), .A2(n2882), .B1(n985), .B2(n3084), .ZN(n2747)
         );
  OAI22_X1 U1076 ( .A1(n3081), .A2(n2883), .B1(n997), .B2(n2343), .ZN(n2736)
         );
  OAI22_X1 U1077 ( .A1(n3081), .A2(n2884), .B1(n992), .B2(n2343), .ZN(n2646)
         );
  OAI22_X1 U1078 ( .A1(n3079), .A2(n2885), .B1(n988), .B2(n3084), .ZN(n2681)
         );
  NAND4_X1 U1079 ( .A1(n2807), .A2(n2808), .A3(n2809), .A4(n2810), .ZN(N103)
         );
  AOI221_X1 U1080 ( .B1(n642), .B2(n3057), .C1(n140), .C2(n3067), .A(n2813), 
        .ZN(n2809) );
  AOI221_X1 U1081 ( .B1(n1891), .B2(n2525), .C1(n646), .C2(n2526), .A(n2814), 
        .ZN(n2808) );
  NAND4_X1 U1082 ( .A1(n2518), .A2(n2519), .A3(n2520), .A4(n2521), .ZN(N99) );
  AOI221_X1 U1083 ( .B1(n194), .B2(n3056), .C1(n143), .C2(n3073), .A(n2524), 
        .ZN(n2520) );
  AOI221_X1 U1084 ( .B1(n1941), .B2(n2525), .C1(n198), .C2(n2526), .A(n2527), 
        .ZN(n2519) );
  NAND4_X1 U1085 ( .A1(n2564), .A2(n2565), .A3(n2566), .A4(n2567), .ZN(N95) );
  AOI221_X1 U1086 ( .B1(n258), .B2(n3052), .C1(n43), .C2(n3069), .A(n2570), 
        .ZN(n2566) );
  AOI221_X1 U1087 ( .B1(n1943), .B2(n2525), .C1(n262), .C2(n2526), .A(n2571), 
        .ZN(n2565) );
  NAND4_X1 U1088 ( .A1(n2608), .A2(n2609), .A3(n2610), .A4(n2611), .ZN(N91) );
  AOI221_X1 U1089 ( .B1(n322), .B2(n3055), .C1(n92), .C2(n3065), .A(n2614), 
        .ZN(n2610) );
  AOI221_X1 U1090 ( .B1(n1539), .B2(n2525), .C1(n326), .C2(n2526), .A(n2615), 
        .ZN(n2609) );
  NAND4_X1 U1091 ( .A1(n2719), .A2(n2720), .A3(n2721), .A4(n2722), .ZN(N111)
         );
  AOI221_X1 U1092 ( .B1(n514), .B2(n3057), .C1(n5), .C2(n3075), .A(n2725), 
        .ZN(n2721) );
  AOI221_X1 U1093 ( .B1(n1475), .B2(n2525), .C1(n518), .C2(n2526), .A(n2726), 
        .ZN(n2720) );
  NAND4_X1 U1094 ( .A1(n2763), .A2(n2764), .A3(n2765), .A4(n2766), .ZN(N107)
         );
  AOI221_X1 U1095 ( .B1(n578), .B2(n3061), .C1(n59), .C2(n3071), .A(n2769), 
        .ZN(n2765) );
  AOI221_X1 U1096 ( .B1(n1478), .B2(n2525), .C1(n582), .C2(n2526), .A(n2770), 
        .ZN(n2764) );
  OAI22_X1 U1097 ( .A1(n831), .A2(n3027), .B1(n863), .B2(n2355), .ZN(n2636) );
  OAI22_X1 U1098 ( .A1(n822), .A2(n3028), .B1(n854), .B2(n3037), .ZN(n2814) );
  OAI22_X1 U1099 ( .A1(n3028), .A2(n2886), .B1(n872), .B2(n3038), .ZN(n2803)
         );
  OAI22_X1 U1100 ( .A1(n823), .A2(n3029), .B1(n855), .B2(n3039), .ZN(n2792) );
  OAI22_X1 U1101 ( .A1(n839), .A2(n3031), .B1(n871), .B2(n3040), .ZN(n2781) );
  OAI22_X1 U1102 ( .A1(n820), .A2(n3030), .B1(n852), .B2(n3043), .ZN(n2527) );
  OAI22_X1 U1103 ( .A1(n842), .A2(n3027), .B1(n874), .B2(n3034), .ZN(n2856) );
  OAI22_X1 U1104 ( .A1(n3032), .A2(n2887), .B1(n853), .B2(n3035), .ZN(n2836)
         );
  OAI22_X1 U1105 ( .A1(n3031), .A2(n2888), .B1(n873), .B2(n3036), .ZN(n2825)
         );
  OAI22_X1 U1106 ( .A1(n818), .A2(n3030), .B1(n850), .B2(n3039), .ZN(n2571) );
  OAI22_X1 U1107 ( .A1(n844), .A2(n3031), .B1(n876), .B2(n3040), .ZN(n2560) );
  OAI22_X1 U1108 ( .A1(n819), .A2(n3032), .B1(n851), .B2(n3041), .ZN(n2549) );
  OAI22_X1 U1109 ( .A1(n843), .A2(n3028), .B1(n875), .B2(n3042), .ZN(n2538) );
  OAI22_X1 U1110 ( .A1(n816), .A2(n3029), .B1(n848), .B2(n3035), .ZN(n2615) );
  OAI22_X1 U1111 ( .A1(n846), .A2(n3029), .B1(n878), .B2(n3036), .ZN(n2604) );
  OAI22_X1 U1112 ( .A1(n3032), .A2(n2889), .B1(n849), .B2(n3037), .ZN(n2593)
         );
  OAI22_X1 U1113 ( .A1(n3027), .A2(n2890), .B1(n877), .B2(n3038), .ZN(n2582)
         );
  OAI22_X1 U1114 ( .A1(n826), .A2(n3032), .B1(n858), .B2(n3045), .ZN(n2726) );
  OAI22_X1 U1115 ( .A1(n836), .A2(n3032), .B1(n868), .B2(n3046), .ZN(n2715) );
  OAI22_X1 U1116 ( .A1(n827), .A2(n3028), .B1(n859), .B2(n3048), .ZN(n2704) );
  OAI22_X1 U1117 ( .A1(n835), .A2(n3028), .B1(n867), .B2(n3045), .ZN(n2693) );
  OAI22_X1 U1118 ( .A1(n824), .A2(n3027), .B1(n856), .B2(n3041), .ZN(n2770) );
  OAI22_X1 U1119 ( .A1(n838), .A2(n3027), .B1(n870), .B2(n3042), .ZN(n2759) );
  OAI22_X1 U1120 ( .A1(n825), .A2(n3030), .B1(n857), .B2(n3043), .ZN(n2748) );
  OAI22_X1 U1121 ( .A1(n837), .A2(n3031), .B1(n869), .B2(n3044), .ZN(n2737) );
  OAI22_X1 U1122 ( .A1(n3031), .A2(n2891), .B1(n879), .B2(n3034), .ZN(n2626)
         );
  OAI22_X1 U1123 ( .A1(n832), .A2(n3029), .B1(n864), .B2(n3048), .ZN(n2647) );
  OAI22_X1 U1124 ( .A1(n828), .A2(n3027), .B1(n860), .B2(n3044), .ZN(n2682) );
  OAI22_X1 U1125 ( .A1(n958), .A2(n3010), .B1(n894), .B2(n3002), .ZN(n2656) );
  OAI22_X1 U1126 ( .A1(n797), .A2(n3020), .B1(n829), .B2(n3030), .ZN(n2669) );
  OAI22_X1 U1127 ( .A1(n927), .A2(n2349), .B1(n799), .B2(n3023), .ZN(n2639) );
  OAI22_X1 U1128 ( .A1(n919), .A2(n2349), .B1(n791), .B2(n3021), .ZN(n2795) );
  OAI22_X1 U1129 ( .A1(n916), .A2(n3017), .B1(n788), .B2(n3022), .ZN(n2530) );
  OAI22_X1 U1130 ( .A1(n914), .A2(n2349), .B1(n786), .B2(n3024), .ZN(n2574) );
  OAI22_X1 U1131 ( .A1(n915), .A2(n3018), .B1(n787), .B2(n3021), .ZN(n2552) );
  OAI22_X1 U1132 ( .A1(n939), .A2(n2349), .B1(n811), .B2(n3022), .ZN(n2541) );
  OAI22_X1 U1133 ( .A1(n912), .A2(n3018), .B1(n784), .B2(n3024), .ZN(n2618) );
  OAI22_X1 U1134 ( .A1(n913), .A2(n3017), .B1(n785), .B2(n3021), .ZN(n2596) );
  OAI22_X1 U1135 ( .A1(n941), .A2(n3018), .B1(n813), .B2(n3022), .ZN(n2585) );
  OAI22_X1 U1136 ( .A1(n920), .A2(n3018), .B1(n792), .B2(n3024), .ZN(n2773) );
  NAND4_X1 U1137 ( .A1(n2640), .A2(n2641), .A3(n2642), .A4(n2643), .ZN(N120)
         );
  AOI221_X1 U1138 ( .B1(n370), .B2(n3053), .C1(n138), .C2(n3078), .A(n2646), 
        .ZN(n2642) );
  AOI221_X1 U1139 ( .B1(n1795), .B2(n2525), .C1(n374), .C2(n2526), .A(n2647), 
        .ZN(n2641) );
  INV_X1 U1140 ( .A(n2648), .ZN(n2640) );
  NAND2_X1 U1141 ( .A1(n2657), .A2(n2658), .ZN(N118) );
  AOI221_X1 U1142 ( .B1(n1958), .B2(n2659), .C1(n1918), .C2(n3077), .A(n2660), 
        .ZN(n2658) );
  AOI221_X1 U1143 ( .B1(n1961), .B2(n2525), .C1(n2661), .C2(n2955), .A(n2663), 
        .ZN(n2657) );
  NAND4_X1 U1144 ( .A1(n2619), .A2(n2620), .A3(n2621), .A4(n2622), .ZN(N90) );
  AOI221_X1 U1145 ( .B1(n338), .B2(n3054), .C1(n96), .C2(n3064), .A(n2625), 
        .ZN(n2621) );
  AOI221_X1 U1146 ( .B1(n1570), .B2(n2525), .C1(n342), .C2(n2526), .A(n2626), 
        .ZN(n2620) );
  INV_X1 U1147 ( .A(n2627), .ZN(n2619) );
  NAND4_X1 U1148 ( .A1(n2675), .A2(n2676), .A3(n2677), .A4(n2678), .ZN(N115)
         );
  AOI221_X1 U1149 ( .B1(n450), .B2(n3062), .C1(n3), .C2(n3074), .A(n2681), 
        .ZN(n2677) );
  AOI221_X1 U1150 ( .B1(n1886), .B2(n2525), .C1(n454), .C2(n2526), .A(n2682), 
        .ZN(n2676) );
  NAND4_X1 U1151 ( .A1(n2796), .A2(n2797), .A3(n2798), .A4(n2799), .ZN(N104)
         );
  AOI221_X1 U1152 ( .B1(n626), .B2(n3058), .C1(n7), .C2(n3068), .A(n2802), 
        .ZN(n2798) );
  AOI221_X1 U1153 ( .B1(n1890), .B2(n2525), .C1(n630), .C2(n2526), .A(n2803), 
        .ZN(n2797) );
  INV_X1 U1154 ( .A(n2804), .ZN(n2796) );
  NAND4_X1 U1155 ( .A1(n2785), .A2(n2786), .A3(n2787), .A4(n2788), .ZN(N105)
         );
  AOI221_X1 U1156 ( .B1(n610), .B2(n3052), .C1(n61), .C2(n3069), .A(n2791), 
        .ZN(n2787) );
  AOI221_X1 U1157 ( .B1(n1889), .B2(n2525), .C1(n614), .C2(n2526), .A(n2792), 
        .ZN(n2786) );
  AOI221_X1 U1158 ( .B1(n613), .B2(n3085), .C1(n2504), .C2(n2933), .A(n2790), 
        .ZN(n2788) );
  NAND4_X1 U1159 ( .A1(n2774), .A2(n2775), .A3(n2776), .A4(n2777), .ZN(N106)
         );
  AOI221_X1 U1160 ( .B1(n594), .B2(n3060), .C1(n6), .C2(n3070), .A(n2780), 
        .ZN(n2776) );
  AOI221_X1 U1161 ( .B1(n1888), .B2(n2525), .C1(n598), .C2(n2526), .A(n2781), 
        .ZN(n2775) );
  INV_X1 U1162 ( .A(n2782), .ZN(n2774) );
  NAND4_X1 U1163 ( .A1(n2840), .A2(n2841), .A3(n2842), .A4(n2843), .ZN(N100)
         );
  AOI221_X1 U1164 ( .B1(n690), .B2(n3054), .C1(n142), .C2(n3064), .A(n2852), 
        .ZN(n2842) );
  AOI221_X1 U1165 ( .B1(n1893), .B2(n2525), .C1(n700), .C2(n2526), .A(n2856), 
        .ZN(n2841) );
  AOI221_X1 U1166 ( .B1(n699), .B2(n3086), .C1(n2504), .C2(n2934), .A(n2845), 
        .ZN(n2843) );
  NAND4_X1 U1167 ( .A1(n2829), .A2(n2830), .A3(n2831), .A4(n2832), .ZN(N101)
         );
  AOI221_X1 U1168 ( .B1(n674), .B2(n3055), .C1(n141), .C2(n3065), .A(n2835), 
        .ZN(n2831) );
  AOI221_X1 U1169 ( .B1(n1940), .B2(n2525), .C1(n678), .C2(n2526), .A(n2836), 
        .ZN(n2830) );
  AOI221_X1 U1170 ( .B1(n677), .B2(n2081), .C1(n2504), .C2(n2935), .A(n2834), 
        .ZN(n2832) );
  NAND4_X1 U1171 ( .A1(n2818), .A2(n2819), .A3(n2820), .A4(n2821), .ZN(N102)
         );
  AOI221_X1 U1172 ( .B1(n658), .B2(n3056), .C1(n9), .C2(n3066), .A(n2824), 
        .ZN(n2820) );
  AOI221_X1 U1173 ( .B1(n1892), .B2(n2525), .C1(n662), .C2(n2526), .A(n2825), 
        .ZN(n2819) );
  AOI221_X1 U1174 ( .B1(n661), .B2(n3085), .C1(n2504), .C2(n2936), .A(n2823), 
        .ZN(n2821) );
  NAND4_X1 U1175 ( .A1(n2553), .A2(n2554), .A3(n2555), .A4(n2556), .ZN(N96) );
  AOI221_X1 U1176 ( .B1(n242), .B2(n3053), .C1(n145), .C2(n3070), .A(n2559), 
        .ZN(n2555) );
  AOI221_X1 U1177 ( .B1(n1506), .B2(n2525), .C1(n246), .C2(n2526), .A(n2560), 
        .ZN(n2554) );
  AOI221_X1 U1178 ( .B1(n245), .B2(n3086), .C1(n2504), .C2(n2937), .A(n2558), 
        .ZN(n2556) );
  NAND4_X1 U1179 ( .A1(n2542), .A2(n2543), .A3(n2544), .A4(n2545), .ZN(N97) );
  AOI221_X1 U1180 ( .B1(n226), .B2(n3054), .C1(n42), .C2(n3071), .A(n2548), 
        .ZN(n2544) );
  AOI221_X1 U1181 ( .B1(n1942), .B2(n2525), .C1(n230), .C2(n2526), .A(n2549), 
        .ZN(n2543) );
  AOI221_X1 U1182 ( .B1(n229), .B2(n2081), .C1(n2504), .C2(n2938), .A(n2547), 
        .ZN(n2545) );
  NAND4_X1 U1183 ( .A1(n2531), .A2(n2532), .A3(n2533), .A4(n2534), .ZN(N98) );
  AOI221_X1 U1184 ( .B1(n210), .B2(n3055), .C1(n144), .C2(n3072), .A(n2537), 
        .ZN(n2533) );
  AOI221_X1 U1185 ( .B1(n1894), .B2(n2525), .C1(n214), .C2(n2526), .A(n2538), 
        .ZN(n2532) );
  AOI221_X1 U1186 ( .B1(n213), .B2(n3085), .C1(n2504), .C2(n2939), .A(n2536), 
        .ZN(n2534) );
  NAND4_X1 U1187 ( .A1(n2597), .A2(n2598), .A3(n2599), .A4(n2600), .ZN(N92) );
  AOI221_X1 U1188 ( .B1(n306), .B2(n3056), .C1(n89), .C2(n3066), .A(n2603), 
        .ZN(n2599) );
  AOI221_X1 U1189 ( .B1(n1538), .B2(n2525), .C1(n310), .C2(n2526), .A(n2604), 
        .ZN(n2598) );
  INV_X1 U1190 ( .A(n2605), .ZN(n2597) );
  NAND4_X1 U1191 ( .A1(n2586), .A2(n2587), .A3(n2588), .A4(n2589), .ZN(N93) );
  AOI221_X1 U1192 ( .B1(n290), .B2(n3057), .C1(n44), .C2(n3067), .A(n2592), 
        .ZN(n2588) );
  AOI221_X1 U1193 ( .B1(n1858), .B2(n2525), .C1(n294), .C2(n2526), .A(n2593), 
        .ZN(n2587) );
  AOI221_X1 U1194 ( .B1(n293), .B2(n3086), .C1(n2504), .C2(n2940), .A(n2591), 
        .ZN(n2589) );
  NAND4_X1 U1195 ( .A1(n2575), .A2(n2576), .A3(n2577), .A4(n2578), .ZN(N94) );
  AOI221_X1 U1196 ( .B1(n274), .B2(n3058), .C1(n88), .C2(n3068), .A(n2581), 
        .ZN(n2577) );
  AOI221_X1 U1197 ( .B1(n1831), .B2(n2525), .C1(n278), .C2(n2526), .A(n2582), 
        .ZN(n2576) );
  AOI221_X1 U1198 ( .B1(n277), .B2(n2081), .C1(n2504), .C2(n2941), .A(n2580), 
        .ZN(n2578) );
  NAND4_X1 U1199 ( .A1(n2708), .A2(n2709), .A3(n2710), .A4(n2711), .ZN(N112)
         );
  AOI221_X1 U1200 ( .B1(n498), .B2(n3059), .C1(n52), .C2(n3076), .A(n2714), 
        .ZN(n2710) );
  AOI221_X1 U1201 ( .B1(n1446), .B2(n2525), .C1(n502), .C2(n2526), .A(n2715), 
        .ZN(n2709) );
  AOI221_X1 U1202 ( .B1(n501), .B2(n3086), .C1(n2504), .C2(n2942), .A(n2713), 
        .ZN(n2711) );
  NAND4_X1 U1203 ( .A1(n2697), .A2(n2698), .A3(n2699), .A4(n2700), .ZN(N113)
         );
  AOI221_X1 U1204 ( .B1(n482), .B2(n3060), .C1(n4), .C2(n3078), .A(n2703), 
        .ZN(n2699) );
  AOI221_X1 U1205 ( .B1(n1411), .B2(n2525), .C1(n486), .C2(n2526), .A(n2704), 
        .ZN(n2698) );
  AOI221_X1 U1206 ( .B1(n485), .B2(n2081), .C1(n2504), .C2(n2943), .A(n2702), 
        .ZN(n2700) );
  NAND4_X1 U1207 ( .A1(n2686), .A2(n2687), .A3(n2688), .A4(n2689), .ZN(N114)
         );
  AOI221_X1 U1208 ( .B1(n466), .B2(n3061), .C1(n139), .C2(n3075), .A(n2692), 
        .ZN(n2688) );
  AOI221_X1 U1209 ( .B1(n1799), .B2(n2525), .C1(n470), .C2(n2526), .A(n2693), 
        .ZN(n2687) );
  AOI221_X1 U1210 ( .B1(n469), .B2(n3085), .C1(n2504), .C2(n2944), .A(n2691), 
        .ZN(n2689) );
  NAND4_X1 U1211 ( .A1(n2752), .A2(n2753), .A3(n2754), .A4(n2755), .ZN(N108)
         );
  AOI221_X1 U1212 ( .B1(n562), .B2(n3062), .C1(n58), .C2(n3072), .A(n2758), 
        .ZN(n2754) );
  AOI221_X1 U1213 ( .B1(n1887), .B2(n2525), .C1(n566), .C2(n2526), .A(n2759), 
        .ZN(n2753) );
  INV_X1 U1214 ( .A(n2760), .ZN(n2752) );
  NAND4_X1 U1215 ( .A1(n2741), .A2(n2742), .A3(n2743), .A4(n2744), .ZN(N109)
         );
  AOI221_X1 U1216 ( .B1(n546), .B2(n3051), .C1(n56), .C2(n3073), .A(n2747), 
        .ZN(n2743) );
  AOI221_X1 U1217 ( .B1(n1830), .B2(n2525), .C1(n550), .C2(n2526), .A(n2748), 
        .ZN(n2742) );
  INV_X1 U1218 ( .A(n2749), .ZN(n2741) );
  NAND4_X1 U1219 ( .A1(n2730), .A2(n2731), .A3(n2732), .A4(n2733), .ZN(N110)
         );
  AOI221_X1 U1220 ( .B1(n530), .B2(n3052), .C1(n55), .C2(n3074), .A(n2736), 
        .ZN(n2732) );
  AOI221_X1 U1221 ( .B1(n1826), .B2(n2525), .C1(n534), .C2(n2526), .A(n2737), 
        .ZN(n2731) );
  AOI221_X1 U1222 ( .B1(n533), .B2(n2081), .C1(n2504), .C2(n2945), .A(n2735), 
        .ZN(n2733) );
  INV_X1 U1223 ( .A(CURR_PC[2]), .ZN(n2862) );
  INV_X1 U1224 ( .A(CURR_PC[4]), .ZN(n2855) );
  INV_X1 U1225 ( .A(CURR_PC[5]), .ZN(n2860) );
  INV_X1 U1226 ( .A(CURR_PC[3]), .ZN(n2861) );
  NAND2_X1 U1227 ( .A1(n2651), .A2(n2652), .ZN(N119) );
  AOI221_X1 U1228 ( .B1(n390), .B2(n2526), .C1(n2510), .C2(n2956), .A(n2656), 
        .ZN(n2651) );
  AOI221_X1 U1229 ( .B1(n2504), .B2(n2958), .C1(n1960), .C2(n2525), .A(n2654), 
        .ZN(n2652) );
  NAND2_X1 U1230 ( .A1(n2664), .A2(n2665), .ZN(N117) );
  AOI221_X1 U1231 ( .B1(n418), .B2(n3051), .C1(n2509), .C2(n2957), .A(n2669), 
        .ZN(n2664) );
  AOI221_X1 U1232 ( .B1(n2504), .B2(n2959), .C1(n1959), .C2(n2659), .A(n2667), 
        .ZN(n2665) );
  OR3_X1 U1233 ( .A1(n2670), .A2(n2671), .A3(n2672), .ZN(N116) );
  OAI22_X1 U1234 ( .A1(n3025), .A2(n802), .B1(n3017), .B2(n930), .ZN(n2671) );
  OAI22_X1 U1235 ( .A1(n3004), .A2(n898), .B1(n3011), .B2(n962), .ZN(n2670) );
  NAND4_X1 U1236 ( .A1(n2630), .A2(n2631), .A3(n2632), .A4(n2633), .ZN(N121)
         );
  AOI221_X1 U1237 ( .B1(n354), .B2(n3053), .C1(n137), .C2(n3077), .A(n2635), 
        .ZN(n2632) );
  AOI221_X1 U1238 ( .B1(n1885), .B2(n2525), .C1(n358), .C2(n2526), .A(n2636), 
        .ZN(n2631) );
  OAI221_X1 U1239 ( .B1(n3007), .B2(n904), .C1(n3013), .C2(n968), .A(n2805), 
        .ZN(n2804) );
  INV_X1 U1240 ( .A(n2806), .ZN(n2805) );
  OAI22_X1 U1241 ( .A1(n936), .A2(n3018), .B1(n808), .B2(n3025), .ZN(n2806) );
  OAI221_X1 U1242 ( .B1(n3007), .B2(n896), .C1(n3012), .C2(n960), .A(n2649), 
        .ZN(n2648) );
  INV_X1 U1243 ( .A(n2650), .ZN(n2649) );
  OAI22_X1 U1244 ( .A1(n928), .A2(n3018), .B1(n800), .B2(n3021), .ZN(n2650) );
  INV_X1 U1245 ( .A(n2837), .ZN(n2829) );
  OAI221_X1 U1246 ( .B1(n3002), .B2(n885), .C1(n3012), .C2(n949), .A(n2838), 
        .ZN(n2837) );
  INV_X1 U1247 ( .A(n2839), .ZN(n2838) );
  OAI22_X1 U1248 ( .A1(n917), .A2(n3018), .B1(n789), .B2(n3021), .ZN(n2839) );
  INV_X1 U1249 ( .A(n2550), .ZN(n2542) );
  OAI221_X1 U1250 ( .B1(n3006), .B2(n883), .C1(n3010), .C2(n947), .A(n2551), 
        .ZN(n2550) );
  INV_X1 U1251 ( .A(n2552), .ZN(n2551) );
  INV_X1 U1252 ( .A(n2616), .ZN(n2608) );
  OAI221_X1 U1253 ( .B1(n3007), .B2(n880), .C1(n3014), .C2(n944), .A(n2617), 
        .ZN(n2616) );
  INV_X1 U1254 ( .A(n2618), .ZN(n2617) );
  INV_X1 U1255 ( .A(n2583), .ZN(n2575) );
  OAI221_X1 U1256 ( .B1(n3006), .B2(n909), .C1(n3015), .C2(n973), .A(n2584), 
        .ZN(n2583) );
  INV_X1 U1257 ( .A(n2585), .ZN(n2584) );
  INV_X1 U1258 ( .A(n2705), .ZN(n2697) );
  OAI221_X1 U1259 ( .B1(n3002), .B2(n891), .C1(n3012), .C2(n955), .A(n2706), 
        .ZN(n2705) );
  INV_X1 U1260 ( .A(n2707), .ZN(n2706) );
  OAI22_X1 U1261 ( .A1(n923), .A2(n3018), .B1(n795), .B2(n3021), .ZN(n2707) );
  INV_X1 U1262 ( .A(n2771), .ZN(n2763) );
  OAI221_X1 U1263 ( .B1(n3005), .B2(n888), .C1(n3014), .C2(n952), .A(n2772), 
        .ZN(n2771) );
  INV_X1 U1264 ( .A(n2773), .ZN(n2772) );
  OAI221_X1 U1265 ( .B1(n3004), .B2(n903), .C1(n3015), .C2(n967), .A(n2783), 
        .ZN(n2782) );
  INV_X1 U1266 ( .A(n2784), .ZN(n2783) );
  OAI22_X1 U1267 ( .A1(n935), .A2(n3017), .B1(n807), .B2(n3023), .ZN(n2784) );
  OAI221_X1 U1268 ( .B1(n3004), .B2(n889), .C1(n3012), .C2(n953), .A(n2750), 
        .ZN(n2749) );
  INV_X1 U1269 ( .A(n2751), .ZN(n2750) );
  OAI22_X1 U1270 ( .A1(n921), .A2(n3017), .B1(n793), .B2(n3025), .ZN(n2751) );
  OAI221_X1 U1271 ( .B1(n3007), .B2(n911), .C1(n3013), .C2(n975), .A(n2628), 
        .ZN(n2627) );
  INV_X1 U1272 ( .A(n2629), .ZN(n2628) );
  OAI22_X1 U1273 ( .A1(n943), .A2(n3017), .B1(n815), .B2(n3023), .ZN(n2629) );
  INV_X1 U1274 ( .A(n2815), .ZN(n2807) );
  OAI221_X1 U1275 ( .B1(n3003), .B2(n886), .C1(n3014), .C2(n950), .A(n2816), 
        .ZN(n2815) );
  INV_X1 U1276 ( .A(n2817), .ZN(n2816) );
  OAI22_X1 U1277 ( .A1(n918), .A2(n3017), .B1(n790), .B2(n3024), .ZN(n2817) );
  INV_X1 U1278 ( .A(n2528), .ZN(n2518) );
  OAI221_X1 U1279 ( .B1(n3007), .B2(n884), .C1(n3011), .C2(n948), .A(n2529), 
        .ZN(n2528) );
  INV_X1 U1280 ( .A(n2530), .ZN(n2529) );
  INV_X1 U1281 ( .A(n2594), .ZN(n2586) );
  OAI221_X1 U1282 ( .B1(n3004), .B2(n881), .C1(n3016), .C2(n945), .A(n2595), 
        .ZN(n2594) );
  INV_X1 U1283 ( .A(n2596), .ZN(n2595) );
  INV_X1 U1284 ( .A(n2637), .ZN(n2630) );
  OAI221_X1 U1285 ( .B1(n2352), .B2(n895), .C1(n2346), .C2(n959), .A(n2638), 
        .ZN(n2637) );
  INV_X1 U1286 ( .A(n2639), .ZN(n2638) );
  INV_X1 U1287 ( .A(n2857), .ZN(n2840) );
  OAI221_X1 U1288 ( .B1(n3003), .B2(n906), .C1(n3011), .C2(n970), .A(n2858), 
        .ZN(n2857) );
  INV_X1 U1289 ( .A(n2859), .ZN(n2858) );
  OAI22_X1 U1290 ( .A1(n938), .A2(n3017), .B1(n810), .B2(n3020), .ZN(n2859) );
  INV_X1 U1291 ( .A(n2561), .ZN(n2553) );
  OAI221_X1 U1292 ( .B1(n3003), .B2(n908), .C1(n3011), .C2(n972), .A(n2562), 
        .ZN(n2561) );
  INV_X1 U1293 ( .A(n2563), .ZN(n2562) );
  OAI22_X1 U1294 ( .A1(n940), .A2(n3017), .B1(n812), .B2(n3020), .ZN(n2563) );
  INV_X1 U1295 ( .A(n2716), .ZN(n2708) );
  OAI221_X1 U1296 ( .B1(n3006), .B2(n900), .C1(n3015), .C2(n964), .A(n2717), 
        .ZN(n2716) );
  INV_X1 U1297 ( .A(n2718), .ZN(n2717) );
  OAI22_X1 U1298 ( .A1(n932), .A2(n3017), .B1(n804), .B2(n3020), .ZN(n2718) );
  INV_X1 U1299 ( .A(n2738), .ZN(n2730) );
  OAI221_X1 U1300 ( .B1(n3005), .B2(n901), .C1(n3012), .C2(n965), .A(n2739), 
        .ZN(n2738) );
  INV_X1 U1301 ( .A(n2740), .ZN(n2739) );
  OAI22_X1 U1302 ( .A1(n933), .A2(n3018), .B1(n805), .B2(n3020), .ZN(n2740) );
  INV_X1 U1303 ( .A(n2683), .ZN(n2675) );
  OAI221_X1 U1304 ( .B1(n3002), .B2(n892), .C1(n3012), .C2(n956), .A(n2684), 
        .ZN(n2683) );
  INV_X1 U1305 ( .A(n2685), .ZN(n2684) );
  OAI22_X1 U1306 ( .A1(n924), .A2(n3017), .B1(n796), .B2(n3020), .ZN(n2685) );
  OAI221_X1 U1307 ( .B1(n3005), .B2(n910), .C1(n3016), .C2(n974), .A(n2606), 
        .ZN(n2605) );
  INV_X1 U1308 ( .A(n2607), .ZN(n2606) );
  OAI22_X1 U1309 ( .A1(n942), .A2(n2349), .B1(n814), .B2(n3025), .ZN(n2607) );
  OAI221_X1 U1310 ( .B1(n3005), .B2(n902), .C1(n3010), .C2(n966), .A(n2761), 
        .ZN(n2760) );
  INV_X1 U1311 ( .A(n2762), .ZN(n2761) );
  OAI22_X1 U1312 ( .A1(n934), .A2(n2349), .B1(n806), .B2(n3025), .ZN(n2762) );
  INV_X1 U1313 ( .A(n2793), .ZN(n2785) );
  OAI221_X1 U1314 ( .B1(n3004), .B2(n887), .C1(n3016), .C2(n951), .A(n2794), 
        .ZN(n2793) );
  INV_X1 U1315 ( .A(n2795), .ZN(n2794) );
  INV_X1 U1316 ( .A(n2826), .ZN(n2818) );
  OAI221_X1 U1317 ( .B1(n3002), .B2(n905), .C1(n3013), .C2(n969), .A(n2827), 
        .ZN(n2826) );
  INV_X1 U1318 ( .A(n2828), .ZN(n2827) );
  OAI22_X1 U1319 ( .A1(n937), .A2(n2349), .B1(n809), .B2(n3022), .ZN(n2828) );
  INV_X1 U1320 ( .A(n2572), .ZN(n2564) );
  OAI221_X1 U1321 ( .B1(n3006), .B2(n882), .C1(n3016), .C2(n946), .A(n2573), 
        .ZN(n2572) );
  INV_X1 U1322 ( .A(n2574), .ZN(n2573) );
  INV_X1 U1323 ( .A(n2539), .ZN(n2531) );
  OAI221_X1 U1324 ( .B1(n3007), .B2(n907), .C1(n3015), .C2(n971), .A(n2540), 
        .ZN(n2539) );
  INV_X1 U1325 ( .A(n2541), .ZN(n2540) );
  INV_X1 U1326 ( .A(n2727), .ZN(n2719) );
  OAI221_X1 U1327 ( .B1(n3003), .B2(n890), .C1(n3010), .C2(n954), .A(n2728), 
        .ZN(n2727) );
  INV_X1 U1328 ( .A(n2729), .ZN(n2728) );
  OAI22_X1 U1329 ( .A1(n922), .A2(n2349), .B1(n794), .B2(n3022), .ZN(n2729) );
  INV_X1 U1330 ( .A(n2694), .ZN(n2686) );
  OAI221_X1 U1331 ( .B1(n3002), .B2(n899), .C1(n3012), .C2(n963), .A(n2695), 
        .ZN(n2694) );
  INV_X1 U1332 ( .A(n2696), .ZN(n2695) );
  OAI22_X1 U1333 ( .A1(n931), .A2(n2349), .B1(n803), .B2(n3022), .ZN(n2696) );
  OAI221_X1 U1334 ( .B1(n2372), .B2(n770), .C1(n3083), .C2(n994), .A(n2673), 
        .ZN(n2672) );
  INV_X1 U1335 ( .A(n2674), .ZN(n2673) );
  OAI22_X1 U1336 ( .A1(n834), .A2(n3028), .B1(n866), .B2(n3047), .ZN(n2674) );
  NOR3_X1 U1337 ( .A1(n749), .A2(n751), .A3(n747), .ZN(n2423) );
  NOR3_X1 U1338 ( .A1(n749), .A2(n751), .A3(n2421), .ZN(n2422) );
  NOR3_X1 U1339 ( .A1(n747), .A2(n749), .A3(n2946), .ZN(n2417) );
  NOR3_X1 U1340 ( .A1(n2946), .A2(n749), .A3(n2421), .ZN(n2415) );
  INV_X1 U1341 ( .A(CURR_PC[1]), .ZN(n2237) );
  INV_X1 U1342 ( .A(CURR_PC[6]), .ZN(n2243) );
  INV_X1 U1343 ( .A(CURR_PC[9]), .ZN(n2233) );
  INV_X1 U1344 ( .A(CURR_PC[10]), .ZN(n2248) );
  INV_X1 U1345 ( .A(CURR_PC[29]), .ZN(n2213) );
  INV_X1 U1346 ( .A(CURR_PC[30]), .ZN(n2268) );
  INV_X1 U1347 ( .A(CURR_PC[14]), .ZN(n2252) );
  INV_X1 U1348 ( .A(CURR_PC[25]), .ZN(n2217) );
  INV_X1 U1349 ( .A(CURR_PC[7]), .ZN(n2235) );
  INV_X1 U1350 ( .A(CURR_PC[8]), .ZN(n2245) );
  INV_X1 U1351 ( .A(CURR_PC[11]), .ZN(n2231) );
  INV_X1 U1352 ( .A(CURR_PC[12]), .ZN(n2250) );
  INV_X1 U1353 ( .A(CURR_PC[27]), .ZN(n2215) );
  INV_X1 U1354 ( .A(CURR_PC[13]), .ZN(n2229) );
  INV_X1 U1355 ( .A(CURR_PC[15]), .ZN(n2227) );
  INV_X1 U1356 ( .A(CURR_PC[16]), .ZN(n2254) );
  INV_X1 U1357 ( .A(CURR_PC[17]), .ZN(n2225) );
  INV_X1 U1358 ( .A(CURR_PC[19]), .ZN(n2223) );
  INV_X1 U1359 ( .A(CURR_PC[21]), .ZN(n2221) );
  INV_X1 U1360 ( .A(CURR_PC[23]), .ZN(n2219) );
  INV_X1 U1361 ( .A(CURR_PC[18]), .ZN(n2256) );
  INV_X1 U1362 ( .A(CURR_PC[20]), .ZN(n2258) );
  INV_X1 U1363 ( .A(CURR_PC[28]), .ZN(n2266) );
  INV_X1 U1364 ( .A(CURR_PC[22]), .ZN(n2260) );
  INV_X1 U1365 ( .A(CURR_PC[24]), .ZN(n2262) );
  INV_X1 U1366 ( .A(CURR_PC[26]), .ZN(n2264) );
  INV_X1 U1367 ( .A(CURR_PC[31]), .ZN(n2210) );
  INV_X1 U1368 ( .A(CURR_PC[0]), .ZN(n2239) );
  NAND2_X1 U1369 ( .A1(n750), .A2(n2947), .ZN(n2424) );
  NAND2_X1 U1370 ( .A1(n750), .A2(n748), .ZN(n2425) );
  OAI22_X1 U1371 ( .A1(n2427), .A2(n2946), .B1(n751), .B2(n2428), .ZN(n2413)
         );
  AOI221_X1 U1372 ( .B1(n2419), .B2(n2432), .C1(n2420), .C2(n2433), .A(n2434), 
        .ZN(n2427) );
  AOI221_X1 U1373 ( .B1(n2419), .B2(n2429), .C1(n2420), .C2(n2430), .A(n2431), 
        .ZN(n2428) );
  OAI22_X1 U1374 ( .A1(n2435), .A2(n2946), .B1(n751), .B2(n2436), .ZN(n2411)
         );
  AOI221_X1 U1375 ( .B1(n2419), .B2(n2440), .C1(n2420), .C2(n2441), .A(n2442), 
        .ZN(n2435) );
  AOI221_X1 U1376 ( .B1(n2419), .B2(n2437), .C1(n2420), .C2(n2438), .A(n2439), 
        .ZN(n2436) );
  AOI211_X1 U1377 ( .C1(n2420), .C2(n2745), .A(n2448), .B(n2421), .ZN(n2446)
         );
  OAI222_X1 U1378 ( .A1(n734), .A2(n2424), .B1(n732), .B2(n2425), .C1(n736), 
        .C2(n2449), .ZN(n2448) );
  AOI211_X1 U1379 ( .C1(n2420), .C2(n2948), .A(n2456), .B(n2421), .ZN(n2454)
         );
  OAI222_X1 U1380 ( .A1(n744), .A2(n2424), .B1(n746), .B2(n2425), .C1(n742), 
        .C2(n2449), .ZN(n2456) );
  OAI221_X1 U1381 ( .B1(n745), .B2(n2425), .C1(n743), .C2(n2424), .A(n2421), 
        .ZN(n2459) );
  AOI221_X1 U1382 ( .B1(n2419), .B2(n2412), .C1(n2420), .C2(n2734), .A(n2452), 
        .ZN(n2445) );
  OAI221_X1 U1383 ( .B1(n733), .B2(n2425), .C1(n735), .C2(n2424), .A(n2421), 
        .ZN(n2452) );
  OAI22_X1 U1384 ( .A1(n719), .A2(n2424), .B1(n717), .B2(n2425), .ZN(n2431) );
  OAI22_X1 U1385 ( .A1(n729), .A2(n2424), .B1(n731), .B2(n2425), .ZN(n2434) );
  OAI22_X1 U1386 ( .A1(n720), .A2(n2424), .B1(n718), .B2(n2425), .ZN(n2439) );
  OAI22_X1 U1387 ( .A1(n728), .A2(n2424), .B1(n730), .B2(n2425), .ZN(n2442) );
  OAI22_X1 U1388 ( .A1(n732), .A2(n2113), .B1(n733), .B2(n2176), .ZN(n2511) );
  OAI22_X1 U1389 ( .A1(n741), .A2(n3018), .B1(n739), .B2(n3023), .ZN(n2515) );
  AND2_X1 U1390 ( .A1(n2443), .A2(n2444), .ZN(n2406) );
  OAI21_X1 U1391 ( .B1(n2453), .B2(n2454), .A(n751), .ZN(n2443) );
  OAI21_X1 U1392 ( .B1(n2445), .B2(n2446), .A(n2946), .ZN(n2444) );
  AOI221_X1 U1393 ( .B1(n2419), .B2(n2949), .C1(n2420), .C2(n2756), .A(n2459), 
        .ZN(n2453) );
  NAND2_X1 U1394 ( .A1(PRED_TK[30]), .A2(n2462), .ZN(n2996) );
  NAND2_X1 U1395 ( .A1(NEXT_PC[30]), .A2(n3094), .ZN(n2997) );
  NAND2_X1 U1397 ( .A1(NEW_PC[30]), .A2(n3098), .ZN(n2998) );
  AOI222_X1 U1398 ( .A1(PRED_TK[31]), .A2(n3091), .B1(NEXT_PC[31]), .B2(n3095), 
        .C1(NEW_PC[31]), .C2(n3098), .ZN(n2471) );
  NOR2_X1 U1399 ( .A1(N815), .A2(n749), .ZN(MISS_HIT[0]) );
  INV_X1 U1400 ( .A(n2471), .ZN(PRED[31]) );
  INV_X1 U1401 ( .A(n2999), .ZN(n3002) );
  INV_X1 U1402 ( .A(n2999), .ZN(n3003) );
  INV_X1 U1403 ( .A(n3000), .ZN(n3004) );
  INV_X1 U1404 ( .A(n3000), .ZN(n3005) );
  INV_X1 U1405 ( .A(n3001), .ZN(n3006) );
  INV_X1 U1406 ( .A(n3001), .ZN(n3007) );
  INV_X1 U1407 ( .A(n3008), .ZN(n3010) );
  INV_X1 U1408 ( .A(n3009), .ZN(n3011) );
  INV_X1 U1409 ( .A(n3009), .ZN(n3012) );
  INV_X1 U1410 ( .A(n3008), .ZN(n3013) );
  INV_X1 U1411 ( .A(n3008), .ZN(n3014) );
  INV_X1 U1412 ( .A(n3008), .ZN(n3015) );
  INV_X1 U1413 ( .A(n3009), .ZN(n3016) );
  BUF_X1 U1414 ( .A(n3033), .Z(n3034) );
  BUF_X1 U1415 ( .A(n3033), .Z(n3035) );
  BUF_X1 U1416 ( .A(n3033), .Z(n3036) );
  BUF_X1 U1417 ( .A(n3033), .Z(n3037) );
  BUF_X1 U1418 ( .A(n3033), .Z(n3038) );
  BUF_X1 U1419 ( .A(n3033), .Z(n3039) );
  BUF_X1 U1420 ( .A(n3033), .Z(n3040) );
  BUF_X1 U1421 ( .A(n3033), .Z(n3041) );
  BUF_X1 U1422 ( .A(n2355), .Z(n3042) );
  BUF_X1 U1423 ( .A(n2355), .Z(n3043) );
  BUF_X1 U1424 ( .A(n2355), .Z(n3044) );
  BUF_X1 U1425 ( .A(n2355), .Z(n3045) );
  BUF_X1 U1426 ( .A(n2355), .Z(n3046) );
  BUF_X1 U1427 ( .A(n2355), .Z(n3047) );
  BUF_X1 U1428 ( .A(n2355), .Z(n3048) );
  BUF_X1 U1429 ( .A(n3063), .Z(n3064) );
  BUF_X1 U1430 ( .A(n3063), .Z(n3065) );
  BUF_X1 U1431 ( .A(n3063), .Z(n3066) );
  BUF_X1 U1432 ( .A(n3063), .Z(n3067) );
  BUF_X1 U1433 ( .A(n3063), .Z(n3068) );
  BUF_X1 U1434 ( .A(n3063), .Z(n3069) );
  BUF_X1 U1435 ( .A(n3063), .Z(n3070) );
  BUF_X1 U1436 ( .A(n3063), .Z(n3071) );
  BUF_X1 U1437 ( .A(n2145), .Z(n3072) );
  BUF_X1 U1438 ( .A(n2145), .Z(n3073) );
  BUF_X1 U1439 ( .A(n2145), .Z(n3074) );
  BUF_X1 U1440 ( .A(n2145), .Z(n3075) );
  BUF_X1 U1441 ( .A(n2145), .Z(n3076) );
  BUF_X1 U1442 ( .A(n2145), .Z(n3077) );
  BUF_X1 U1443 ( .A(n2145), .Z(n3078) );
  INV_X1 U1444 ( .A(n3103), .ZN(n3098) );
  INV_X1 U1445 ( .A(n3100), .ZN(n3099) );
  INV_X1 U1446 ( .A(n3097), .ZN(n3100) );
  INV_X1 U1447 ( .A(n3100), .ZN(n3101) );
  INV_X1 U1448 ( .A(n3100), .ZN(n3102) );
  INV_X1 U1449 ( .A(n2464), .ZN(n3103) );
  INV_X1 U1450 ( .A(n3103), .ZN(n3104) );
  INV_X1 U1451 ( .A(n3103), .ZN(n3105) );
  INV_X1 U1452 ( .A(n2179), .ZN(n3155) );
  INV_X1 U1453 ( .A(n2179), .ZN(n3156) );
  INV_X1 U1454 ( .A(n2116), .ZN(n3161) );
  INV_X1 U1455 ( .A(n2116), .ZN(n3162) );
  INV_X1 U1456 ( .A(n2053), .ZN(n3167) );
  INV_X1 U1457 ( .A(n2053), .ZN(n3168) );
  BUF_X1 U1458 ( .A(n2246), .Z(n3183) );
  BUF_X1 U1459 ( .A(n2246), .Z(n3184) );
  BUF_X1 U1460 ( .A(n2246), .Z(n3185) );
  BUF_X1 U1461 ( .A(n2246), .Z(n3186) );
  BUF_X1 U1462 ( .A(n2246), .Z(n3187) );
  CLKBUF_X1 U1463 ( .A(n3245), .Z(n3188) );
  CLKBUF_X1 U1464 ( .A(n3245), .Z(n3189) );
  CLKBUF_X1 U1465 ( .A(n3245), .Z(n3190) );
  CLKBUF_X1 U1466 ( .A(n3245), .Z(n3191) );
  CLKBUF_X1 U1467 ( .A(n3244), .Z(n3192) );
  CLKBUF_X1 U1468 ( .A(n3244), .Z(n3193) );
  CLKBUF_X1 U1469 ( .A(n3244), .Z(n3194) );
  CLKBUF_X1 U1470 ( .A(n3244), .Z(n3195) );
  CLKBUF_X1 U1471 ( .A(n3244), .Z(n3196) );
  CLKBUF_X1 U1472 ( .A(n3243), .Z(n3197) );
  CLKBUF_X1 U1473 ( .A(n3243), .Z(n3198) );
  CLKBUF_X1 U1474 ( .A(n3243), .Z(n3199) );
  CLKBUF_X1 U1475 ( .A(n3243), .Z(n3200) );
  CLKBUF_X1 U1476 ( .A(n3243), .Z(n3201) );
  CLKBUF_X1 U1477 ( .A(n3242), .Z(n3202) );
  CLKBUF_X1 U1478 ( .A(n3242), .Z(n3203) );
  CLKBUF_X1 U1479 ( .A(n3242), .Z(n3204) );
  CLKBUF_X1 U1480 ( .A(n3242), .Z(n3205) );
  CLKBUF_X1 U1481 ( .A(n3242), .Z(n3206) );
  CLKBUF_X1 U1482 ( .A(n3241), .Z(n3207) );
  CLKBUF_X1 U1483 ( .A(n3241), .Z(n3208) );
  CLKBUF_X1 U1484 ( .A(n3241), .Z(n3209) );
  CLKBUF_X1 U1485 ( .A(n3241), .Z(n3210) );
  CLKBUF_X1 U1486 ( .A(n3241), .Z(n3211) );
  CLKBUF_X1 U1487 ( .A(n3240), .Z(n3212) );
  CLKBUF_X1 U1488 ( .A(n3240), .Z(n3213) );
  CLKBUF_X1 U1489 ( .A(n3240), .Z(n3214) );
  CLKBUF_X1 U1490 ( .A(n3240), .Z(n3215) );
  CLKBUF_X1 U1491 ( .A(n3240), .Z(n3216) );
  CLKBUF_X1 U1492 ( .A(n3239), .Z(n3217) );
  CLKBUF_X1 U1493 ( .A(n3239), .Z(n3218) );
  CLKBUF_X1 U1494 ( .A(n3239), .Z(n3219) );
  CLKBUF_X1 U1495 ( .A(n3239), .Z(n3220) );
  CLKBUF_X1 U1496 ( .A(n3239), .Z(n3221) );
  CLKBUF_X1 U1497 ( .A(n3238), .Z(n3222) );
  CLKBUF_X1 U1498 ( .A(n3238), .Z(n3223) );
  CLKBUF_X1 U1499 ( .A(n3238), .Z(n3224) );
  CLKBUF_X1 U1500 ( .A(n3238), .Z(n3225) );
  CLKBUF_X1 U1501 ( .A(n3238), .Z(n3226) );
  CLKBUF_X1 U1502 ( .A(n3237), .Z(n3227) );
  CLKBUF_X1 U1503 ( .A(n3237), .Z(n3228) );
  CLKBUF_X1 U1504 ( .A(n3237), .Z(n3229) );
  CLKBUF_X1 U1505 ( .A(n3237), .Z(n3230) );
  CLKBUF_X1 U1506 ( .A(n3237), .Z(n3231) );
  CLKBUF_X1 U1507 ( .A(n3236), .Z(n3232) );
  CLKBUF_X1 U1508 ( .A(n3236), .Z(n3233) );
  CLKBUF_X1 U1509 ( .A(n3236), .Z(n3234) );
  CLKBUF_X1 U1510 ( .A(n3236), .Z(n3235) );
endmodule


module FD_INJ_NB32_0 ( CK, RESET, INJ_ZERO, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   n38, n39, n40, n41, n42, n43, n44;
  wire   [31:0] TMP_D;
  assign n38 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(TMP_D[31]), .CK(CK), .RN(n44), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(TMP_D[30]), .CK(CK), .RN(n44), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(TMP_D[29]), .CK(CK), .RN(n44), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(TMP_D[28]), .CK(CK), .RN(n44), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(TMP_D[27]), .CK(CK), .RN(n44), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(TMP_D[26]), .CK(CK), .RN(n44), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(TMP_D[25]), .CK(CK), .RN(n44), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(TMP_D[24]), .CK(CK), .RN(n44), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(TMP_D[23]), .CK(CK), .RN(n42), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(TMP_D[22]), .CK(CK), .RN(n42), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(TMP_D[21]), .CK(CK), .RN(n42), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(TMP_D[20]), .CK(CK), .RN(n42), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(TMP_D[19]), .CK(CK), .RN(n42), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(TMP_D[18]), .CK(CK), .RN(n42), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(TMP_D[17]), .CK(CK), .RN(n42), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(TMP_D[16]), .CK(CK), .RN(n42), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(TMP_D[15]), .CK(CK), .RN(n42), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(TMP_D[14]), .CK(CK), .RN(n42), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(TMP_D[13]), .CK(CK), .RN(n42), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(TMP_D[12]), .CK(CK), .RN(n42), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(TMP_D[11]), .CK(CK), .RN(n43), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(TMP_D[10]), .CK(CK), .RN(n43), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(TMP_D[9]), .CK(CK), .RN(n43), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(TMP_D[8]), .CK(CK), .RN(n43), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(TMP_D[7]), .CK(CK), .RN(n43), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(TMP_D[6]), .CK(CK), .RN(n43), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(TMP_D[5]), .CK(CK), .RN(n43), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(TMP_D[4]), .CK(CK), .RN(n43), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(TMP_D[3]), .CK(CK), .RN(n43), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(TMP_D[2]), .CK(CK), .RN(n43), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(TMP_D[1]), .CK(CK), .RN(n43), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(TMP_D[0]), .CK(CK), .RN(n43), .Q(Q[0]) );
  BUF_X1 U3 ( .A(n38), .Z(n43) );
  BUF_X1 U4 ( .A(n38), .Z(n42) );
  BUF_X1 U5 ( .A(n38), .Z(n44) );
  AND2_X1 U6 ( .A1(D[3]), .A2(n41), .ZN(TMP_D[3]) );
  AND2_X1 U7 ( .A1(D[4]), .A2(n41), .ZN(TMP_D[4]) );
  AND2_X1 U8 ( .A1(D[6]), .A2(n41), .ZN(TMP_D[6]) );
  AND2_X1 U9 ( .A1(D[7]), .A2(n41), .ZN(TMP_D[7]) );
  AND2_X1 U10 ( .A1(D[10]), .A2(n39), .ZN(TMP_D[10]) );
  AND2_X1 U11 ( .A1(D[11]), .A2(n39), .ZN(TMP_D[11]) );
  AND2_X1 U12 ( .A1(D[14]), .A2(n39), .ZN(TMP_D[14]) );
  AND2_X1 U13 ( .A1(D[5]), .A2(n41), .ZN(TMP_D[5]) );
  AND2_X1 U14 ( .A1(D[8]), .A2(n41), .ZN(TMP_D[8]) );
  AND2_X1 U15 ( .A1(D[15]), .A2(n39), .ZN(TMP_D[15]) );
  AND2_X1 U16 ( .A1(D[16]), .A2(n39), .ZN(TMP_D[16]) );
  AND2_X1 U17 ( .A1(D[17]), .A2(n39), .ZN(TMP_D[17]) );
  AND2_X1 U18 ( .A1(D[18]), .A2(n39), .ZN(TMP_D[18]) );
  AND2_X1 U19 ( .A1(D[22]), .A2(n40), .ZN(TMP_D[22]) );
  AND2_X1 U20 ( .A1(D[23]), .A2(n40), .ZN(TMP_D[23]) );
  AND2_X1 U21 ( .A1(D[12]), .A2(n39), .ZN(TMP_D[12]) );
  AND2_X1 U22 ( .A1(D[13]), .A2(n39), .ZN(TMP_D[13]) );
  AND2_X1 U23 ( .A1(D[19]), .A2(n39), .ZN(TMP_D[19]) );
  AND2_X1 U24 ( .A1(D[21]), .A2(n40), .ZN(TMP_D[21]) );
  AND2_X1 U25 ( .A1(D[24]), .A2(n40), .ZN(TMP_D[24]) );
  AND2_X1 U26 ( .A1(D[25]), .A2(n40), .ZN(TMP_D[25]) );
  AND2_X1 U27 ( .A1(D[26]), .A2(n40), .ZN(TMP_D[26]) );
  AND2_X1 U28 ( .A1(D[29]), .A2(n40), .ZN(TMP_D[29]) );
  AND2_X1 U29 ( .A1(D[28]), .A2(n40), .ZN(TMP_D[28]) );
  AND2_X1 U30 ( .A1(D[20]), .A2(n40), .ZN(TMP_D[20]) );
  AND2_X1 U31 ( .A1(D[27]), .A2(n40), .ZN(TMP_D[27]) );
  AND2_X1 U32 ( .A1(D[30]), .A2(n40), .ZN(TMP_D[30]) );
  AND2_X1 U33 ( .A1(n41), .A2(D[9]), .ZN(TMP_D[9]) );
  AND2_X1 U34 ( .A1(D[31]), .A2(n41), .ZN(TMP_D[31]) );
  AND2_X1 U35 ( .A1(D[2]), .A2(n40), .ZN(TMP_D[2]) );
  AND2_X1 U36 ( .A1(D[0]), .A2(n39), .ZN(TMP_D[0]) );
  AND2_X1 U37 ( .A1(D[1]), .A2(n39), .ZN(TMP_D[1]) );
  CLKBUF_X1 U38 ( .A(INJ_ZERO), .Z(n40) );
  CLKBUF_X1 U39 ( .A(INJ_ZERO), .Z(n41) );
  CLKBUF_X1 U40 ( .A(INJ_ZERO), .Z(n39) );
endmodule


module FD_INJ_NB1_0 ( CK, RESET, INJ_ZERO, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET, INJ_ZERO;
  wire   \TMP_D[0] ;

  DFFR_X1 \Q_reg[0]  ( .D(\TMP_D[0] ), .CK(CK), .RN(RESET), .Q(Q[0]) );
  AND2_X1 U3 ( .A1(INJ_ZERO), .A2(D[0]), .ZN(\TMP_D[0] ) );
endmodule


module FD_NB4_0 ( CK, RESET, D, Q );
  input [3:0] D;
  output [3:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB3_0 ( CK, RESET, D, Q );
  input [2:0] D;
  output [2:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB2_0 ( CK, RESET, D, Q );
  input [1:0] D;
  output [1:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB1_0 ( CK, RESET, D, Q );
  input [0:0] D;
  output [0:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB11_0 ( CK, RESET, D, Q );
  input [10:0] D;
  output [10:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[10]  ( .D(D[10]), .CK(CK), .RN(RESET), .Q(Q[10]) );
  DFFR_X1 \TMP_Q_reg[9]  ( .D(D[9]), .CK(CK), .RN(RESET), .Q(Q[9]) );
  DFFR_X1 \TMP_Q_reg[8]  ( .D(D[8]), .CK(CK), .RN(RESET), .Q(Q[8]) );
  DFFR_X1 \TMP_Q_reg[7]  ( .D(D[7]), .CK(CK), .RN(RESET), .Q(Q[7]) );
  DFFR_X1 \TMP_Q_reg[6]  ( .D(D[6]), .CK(CK), .RN(RESET), .Q(Q[6]) );
  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FD_NB6_0 ( CK, RESET, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET;


  DFFR_X1 \TMP_Q_reg[5]  ( .D(D[5]), .CK(CK), .RN(RESET), .Q(Q[5]) );
  DFFR_X1 \TMP_Q_reg[4]  ( .D(D[4]), .CK(CK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \TMP_Q_reg[3]  ( .D(D[3]), .CK(CK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \TMP_Q_reg[2]  ( .D(D[2]), .CK(CK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \TMP_Q_reg[1]  ( .D(D[1]), .CK(CK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \TMP_Q_reg[0]  ( .D(D[0]), .CK(CK), .RN(RESET), .Q(Q[0]) );
endmodule


module FOREWARD_UNIT_NB32_LS5 ( .INST_EX({\INST_EX[1] , \INST_EX[0] }), 
    .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }), INST_T_EX, Rs_EX, Rt_EX, Rd_MEM, 
        Rd_WB, CTL_MUX1, CTL_MUX2 );
  input [4:0] Rs_EX;
  input [4:0] Rt_EX;
  input [4:0] Rd_MEM;
  input [4:0] Rd_WB;
  output [1:0] CTL_MUX1;
  output [1:0] CTL_MUX2;
  input \INST_EX[1] , \INST_EX[0] , \INST_MEM[1] , \INST_MEM[0] , INST_T_EX;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n57, n58,
         n59;

  XOR2_X1 U39 ( .A(Rt_EX[1]), .B(Rd_MEM[1]), .Z(n25) );
  XOR2_X1 U40 ( .A(Rt_EX[0]), .B(Rd_MEM[0]), .Z(n24) );
  XOR2_X1 U41 ( .A(Rt_EX[4]), .B(Rd_MEM[4]), .Z(n23) );
  XOR2_X1 U42 ( .A(Rs_EX[2]), .B(Rd_WB[2]), .Z(n29) );
  XOR2_X1 U43 ( .A(Rs_EX[1]), .B(Rd_MEM[1]), .Z(n44) );
  XOR2_X1 U44 ( .A(Rs_EX[0]), .B(Rd_MEM[0]), .Z(n43) );
  XOR2_X1 U45 ( .A(Rs_EX[4]), .B(Rd_MEM[4]), .Z(n42) );
  OR3_X1 U2 ( .A1(n28), .A2(n29), .A3(n27), .ZN(n57) );
  NOR2_X1 U3 ( .A1(n26), .A2(n57), .ZN(CTL_MUX1[1]) );
  AND2_X1 U4 ( .A1(n40), .A2(n39), .ZN(n58) );
  NAND2_X1 U5 ( .A1(n30), .A2(n31), .ZN(n38) );
  XNOR2_X1 U6 ( .A(Rs_EX[1]), .B(n31), .ZN(n27) );
  XNOR2_X1 U7 ( .A(Rs_EX[0]), .B(n30), .ZN(n28) );
  INV_X1 U8 ( .A(INST_T_EX), .ZN(n18) );
  NAND4_X1 U9 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .ZN(n10) );
  INV_X1 U10 ( .A(INST_EX[1]), .ZN(n46) );
  OR2_X1 U11 ( .A1(Rd_MEM[0]), .A2(Rd_MEM[1]), .ZN(n48) );
  XNOR2_X1 U12 ( .A(Rd_MEM[3]), .B(Rt_EX[3]), .ZN(n21) );
  XNOR2_X1 U13 ( .A(Rd_WB[1]), .B(Rt_EX[1]), .ZN(n14) );
  XNOR2_X1 U14 ( .A(Rd_WB[2]), .B(Rt_EX[2]), .ZN(n11) );
  XNOR2_X1 U15 ( .A(Rd_WB[4]), .B(Rt_EX[4]), .ZN(n15) );
  AND2_X1 U16 ( .A1(n33), .A2(n32), .ZN(n59) );
  INV_X1 U17 ( .A(Rd_WB[1]), .ZN(n31) );
  OAI22_X1 U18 ( .A1(INST_MEM[0]), .A2(n36), .B1(n37), .B2(n38), .ZN(n35) );
  INV_X1 U19 ( .A(INST_MEM[1]), .ZN(n36) );
  OR3_X1 U20 ( .A1(Rd_MEM[3]), .A2(Rd_MEM[4]), .A3(Rd_MEM[2]), .ZN(n47) );
  NAND3_X1 U21 ( .A1(n34), .A2(n16), .A3(n59), .ZN(n26) );
  NAND3_X1 U22 ( .A1(n20), .A2(n41), .A3(n58), .ZN(n34) );
  XNOR2_X1 U23 ( .A(Rd_WB[4]), .B(Rs_EX[4]), .ZN(n33) );
  XNOR2_X1 U24 ( .A(Rd_MEM[3]), .B(Rs_EX[3]), .ZN(n40) );
  NOR3_X1 U25 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n41) );
  XNOR2_X1 U26 ( .A(Rd_WB[3]), .B(Rt_EX[3]), .ZN(n12) );
  OR3_X1 U27 ( .A1(Rd_WB[3]), .A2(Rd_WB[4]), .A3(Rd_WB[2]), .ZN(n37) );
  XNOR2_X1 U28 ( .A(Rd_WB[3]), .B(Rs_EX[3]), .ZN(n32) );
  INV_X1 U29 ( .A(n34), .ZN(CTL_MUX1[0]) );
  NAND4_X1 U30 ( .A1(n15), .A2(INST_T_EX), .A3(n16), .A4(n17), .ZN(n9) );
  NOR2_X1 U31 ( .A1(n18), .A2(n17), .ZN(CTL_MUX2[0]) );
  NOR2_X1 U32 ( .A1(n9), .A2(n10), .ZN(CTL_MUX2[1]) );
  NOR3_X1 U33 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n22) );
  INV_X1 U34 ( .A(n35), .ZN(n16) );
  XNOR2_X1 U35 ( .A(Rd_WB[0]), .B(Rt_EX[0]), .ZN(n13) );
  INV_X1 U36 ( .A(Rd_WB[0]), .ZN(n30) );
  NAND4_X1 U37 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(n17) );
  OAI22_X1 U38 ( .A1(INST_EX[0]), .A2(n46), .B1(n47), .B2(n48), .ZN(n45) );
  XNOR2_X1 U46 ( .A(Rd_MEM[2]), .B(Rs_EX[2]), .ZN(n39) );
  XNOR2_X1 U47 ( .A(Rd_MEM[2]), .B(Rt_EX[2]), .ZN(n19) );
  INV_X1 U48 ( .A(n45), .ZN(n20) );
endmodule


module WRITE_BACK_UNIT_NB32_LS5 ( MEM_ALU_SEL, DEST_IN, FROM_ALU, FROM_MEM, 
        DATA_OUT, DEST_OUT );
  input [4:0] DEST_IN;
  input [31:0] FROM_ALU;
  input [31:0] FROM_MEM;
  output [31:0] DATA_OUT;
  output [4:0] DEST_OUT;
  input MEM_ALU_SEL;

  assign DEST_OUT[4] = DEST_IN[4];
  assign DEST_OUT[3] = DEST_IN[3];
  assign DEST_OUT[2] = DEST_IN[2];
  assign DEST_OUT[1] = DEST_IN[1];
  assign DEST_OUT[0] = DEST_IN[0];

  MUX21_generic_NB32_1 wb_mux ( .A(FROM_ALU), .B(FROM_MEM), .SEL(MEM_ALU_SEL), 
        .Y(DATA_OUT) );
endmodule


module MEMORY_UNIT_NB32_LS5 ( CLK, RST, DEST_IN, FROM_MEM, FROM_ALU, ALU_OUT, 
        MEM_OUT, DEST_OUT );
  input [4:0] DEST_IN;
  input [31:0] FROM_MEM;
  input [31:0] FROM_ALU;
  output [31:0] ALU_OUT;
  output [31:0] MEM_OUT;
  output [4:0] DEST_OUT;
  input CLK, RST;


  FD_NB32_2 exec_reg ( .CK(CLK), .RESET(RST), .D(FROM_ALU), .Q(ALU_OUT) );
  FD_NB32_1 mem_reg ( .CK(CLK), .RESET(RST), .D(FROM_MEM), .Q(MEM_OUT) );
  FD_NB5_1 dest_reg ( .CK(CLK), .RESET(RST), .D(DEST_IN), .Q(DEST_OUT) );
endmodule


module EXECUTION_UNIT_NB32_LS5 ( FW_MUX1_SEL, FW_MUX2_SEL, FW_EX, FW_MEM, A, B, 
        C, D, DEST_IN, CLK, RST, US, MUX1_SEL, MUX2_SEL, UN_SEL, OP_SEL, 
        US_MEM, TEMP_PC, ALU_OUT, IMM_OUT, DEST_OUT );
  input [1:0] FW_MUX1_SEL;
  input [1:0] FW_MUX2_SEL;
  input [31:0] FW_EX;
  input [31:0] FW_MEM;
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [4:0] DEST_IN;
  input [2:0] UN_SEL;
  input [3:0] OP_SEL;
  output [31:0] TEMP_PC;
  output [31:0] ALU_OUT;
  output [31:0] IMM_OUT;
  output [4:0] DEST_OUT;
  input CLK, RST, US, MUX1_SEL, MUX2_SEL;
  output US_MEM;
  wire   CA_OUT, n1, n2, n3, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49;
  wire   [30:0] TERM1;
  wire   [30:0] TERM2;
  wire   [1:0] MSB;
  wire   [31:0] TERM4;
  wire   [31:0] TERM5;
  wire   [31:0] TERM3;
  wire   [31:0] MUL_OUT;
  wire   [31:0] SHFT_OUT;
  wire   [31:0] COMP_OUT;
  wire   [31:0] LOGIC_OUT;
  wire   [4:0] TMP_DEST_OUT;
  wire   [31:0] MUX2_OUT;
  wire   [31:0] JMP_RET;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  XOR2_X1 U16 ( .A(TERM2[9]), .B(n49), .Z(TERM3[9]) );
  XOR2_X1 U17 ( .A(TERM2[8]), .B(n49), .Z(TERM3[8]) );
  XOR2_X1 U18 ( .A(TERM2[7]), .B(n49), .Z(TERM3[7]) );
  XOR2_X1 U19 ( .A(TERM2[6]), .B(n49), .Z(TERM3[6]) );
  XOR2_X1 U20 ( .A(TERM2[5]), .B(n49), .Z(TERM3[5]) );
  XOR2_X1 U21 ( .A(TERM2[4]), .B(n49), .Z(TERM3[4]) );
  XOR2_X1 U22 ( .A(TERM2[3]), .B(n49), .Z(TERM3[3]) );
  XOR2_X1 U23 ( .A(n49), .B(MSB[0]), .Z(TERM3[31]) );
  XOR2_X1 U24 ( .A(TERM2[30]), .B(n49), .Z(TERM3[30]) );
  XOR2_X1 U25 ( .A(TERM2[2]), .B(n49), .Z(TERM3[2]) );
  XOR2_X1 U26 ( .A(TERM2[29]), .B(n48), .Z(TERM3[29]) );
  XOR2_X1 U27 ( .A(TERM2[28]), .B(n48), .Z(TERM3[28]) );
  XOR2_X1 U28 ( .A(TERM2[27]), .B(n48), .Z(TERM3[27]) );
  XOR2_X1 U29 ( .A(TERM2[26]), .B(n48), .Z(TERM3[26]) );
  XOR2_X1 U30 ( .A(TERM2[25]), .B(n48), .Z(TERM3[25]) );
  XOR2_X1 U31 ( .A(TERM2[24]), .B(n48), .Z(TERM3[24]) );
  XOR2_X1 U32 ( .A(TERM2[23]), .B(n48), .Z(TERM3[23]) );
  XOR2_X1 U33 ( .A(TERM2[22]), .B(n48), .Z(TERM3[22]) );
  XOR2_X1 U34 ( .A(TERM2[21]), .B(n48), .Z(TERM3[21]) );
  XOR2_X1 U35 ( .A(TERM2[20]), .B(n48), .Z(TERM3[20]) );
  XOR2_X1 U36 ( .A(TERM2[1]), .B(n48), .Z(TERM3[1]) );
  XOR2_X1 U37 ( .A(TERM2[19]), .B(n48), .Z(TERM3[19]) );
  XOR2_X1 U38 ( .A(TERM2[18]), .B(n48), .Z(TERM3[18]) );
  XOR2_X1 U39 ( .A(TERM2[17]), .B(n47), .Z(TERM3[17]) );
  XOR2_X1 U40 ( .A(TERM2[16]), .B(n47), .Z(TERM3[16]) );
  XOR2_X1 U41 ( .A(TERM2[15]), .B(n47), .Z(TERM3[15]) );
  XOR2_X1 U42 ( .A(TERM2[14]), .B(n47), .Z(TERM3[14]) );
  XOR2_X1 U43 ( .A(TERM2[13]), .B(n47), .Z(TERM3[13]) );
  XOR2_X1 U44 ( .A(TERM2[12]), .B(n47), .Z(TERM3[12]) );
  XOR2_X1 U45 ( .A(TERM2[11]), .B(n47), .Z(TERM3[11]) );
  XOR2_X1 U46 ( .A(TERM2[10]), .B(n47), .Z(TERM3[10]) );
  MUX21_generic_NB32_3 mux1 ( .A(A), .B(D), .SEL(MUX1_SEL), .Y(TERM4) );
  MUX21_generic_NB32_2 mux2 ( .A(B), .B(C), .SEL(MUX2_SEL), .Y(TERM5) );
  MUX31_generic_NB32_0 fW_mux1 ( .A(TERM4), .B(FW_EX), .C(FW_MEM), .SEL(
        FW_MUX1_SEL), .Y({MSB[1], TERM1[30:16], n21, n20, n19, n18, n17, n16, 
        n15, n14, n13, n12, n11, n10, n9, n3, n2, n1}) );
  MUX31_generic_NB32_1 fw_mux2 ( .A(TERM5), .B(FW_EX), .C(FW_MEM), .SEL(
        FW_MUX2_SEL), .Y({MSB[0], TERM2}) );
  p4addgen_NB32_CW4_0 adder ( .A({MSB[1], TERM1[30:16], n21, n32, n33, n34, 
        n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n1}), .B(TERM3), 
        .Ci(n47), .Co(CA_OUT), .S(TEMP_PC) );
  BOOTHMUL_NB32 multiplier ( .A({n21, n32, n33, n34, n35, n36, n37, n38, n39, 
        n40, n41, n42, n43, n44, n45, n46}), .B({TERM2[15:11], n29, TERM2[9:0]}), .C(MUL_OUT) );
  SHIFTER_NB32_LS5 shift_rot ( .FUNC({OP_SEL[1], n49}), .US(US), .DATA1({
        MSB[1], TERM1[30:16], n21, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
        n41, n42, n43, n44, n45, n46}), .DATA2(TERM2[4:0]), .OUTSHFT(SHFT_OUT)
         );
  COMPARATOR_NB32 comparison ( .AdderRes({TEMP_PC[31:23], n30, n31, 
        TEMP_PC[20:0]}), .MSB(MSB), .CO(CA_OUT), .OP_CODE(OP_SEL[3:1]), .US(US), .SOUT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, COMP_OUT[0]}) );
  LOGIC_NB32 log_un ( .SEL({OP_SEL[3:1], n47}), .A({MSB[1], TERM1[30:16], n21, 
        n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
        n46}), .B({MSB[0], TERM2}), .RES(LOGIC_OUT) );
  FD_NB5_0 destination_register ( .CK(CLK), .RESET(RST), .D(TMP_DEST_OUT), .Q(
        DEST_OUT) );
  FD_NB32_4 output_register ( .CK(CLK), .RESET(RST), .D(MUX2_OUT), .Q(ALU_OUT)
         );
  FD_NB32_3 imm_register ( .CK(CLK), .RESET(RST), .D(B), .Q(IMM_OUT) );
  FD_NB1_1 us_register ( .CK(CLK), .RESET(RST), .D(US), .Q(US_MEM) );
  MUX61_generic_NB32 mux_out ( .A({TEMP_PC[31:23], n30, n31, TEMP_PC[20:0]}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, COMP_OUT[0]}), .C(
        MUL_OUT), .D(SHFT_OUT), .E(LOGIC_OUT), .F(JMP_RET), .SEL(UN_SEL), .Y(
        MUX2_OUT) );
  EXECUTION_UNIT_NB32_LS5_DW01_add_0 add_202 ( .A(D), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(JMP_RET) );
  BUF_X1 U3 ( .A(OP_SEL[0]), .Z(n48) );
  NAND2_X1 U5 ( .A1(TERM2[0]), .A2(n26), .ZN(n27) );
  NAND2_X1 U6 ( .A1(n25), .A2(n48), .ZN(n28) );
  NAND2_X1 U9 ( .A1(n27), .A2(n28), .ZN(TERM3[0]) );
  INV_X1 U10 ( .A(TERM2[0]), .ZN(n25) );
  INV_X1 U11 ( .A(n48), .ZN(n26) );
  BUF_X1 U12 ( .A(n1), .Z(n46) );
  BUF_X2 U13 ( .A(n18), .Z(n34) );
  BUF_X2 U14 ( .A(n10), .Z(n42) );
  BUF_X2 U15 ( .A(n20), .Z(n32) );
  BUF_X2 U47 ( .A(n12), .Z(n40) );
  BUF_X2 U48 ( .A(n3), .Z(n44) );
  BUF_X2 U49 ( .A(n11), .Z(n41) );
  BUF_X1 U50 ( .A(OP_SEL[0]), .Z(n49) );
  BUF_X1 U51 ( .A(OP_SEL[0]), .Z(n47) );
  AND3_X1 U52 ( .A1(OP_SEL[2]), .A2(n49), .A3(n24), .ZN(n23) );
  NOR2_X1 U53 ( .A1(OP_SEL[3]), .A2(OP_SEL[1]), .ZN(n24) );
  OR2_X1 U54 ( .A1(n23), .A2(DEST_IN[0]), .ZN(TMP_DEST_OUT[0]) );
  OR2_X1 U55 ( .A1(n23), .A2(DEST_IN[1]), .ZN(TMP_DEST_OUT[1]) );
  OR2_X1 U56 ( .A1(n23), .A2(DEST_IN[2]), .ZN(TMP_DEST_OUT[2]) );
  OR2_X1 U57 ( .A1(n23), .A2(DEST_IN[3]), .ZN(TMP_DEST_OUT[3]) );
  OR2_X1 U58 ( .A1(n23), .A2(DEST_IN[4]), .ZN(TMP_DEST_OUT[4]) );
  BUF_X1 U59 ( .A(TERM2[10]), .Z(n29) );
  CLKBUF_X1 U60 ( .A(TEMP_PC[22]), .Z(n30) );
  CLKBUF_X1 U61 ( .A(TEMP_PC[21]), .Z(n31) );
  BUF_X4 U62 ( .A(n14), .Z(n38) );
  BUF_X4 U94 ( .A(n16), .Z(n36) );
  BUF_X4 U95 ( .A(n15), .Z(n37) );
  BUF_X4 U96 ( .A(n2), .Z(n45) );
  BUF_X4 U97 ( .A(n17), .Z(n35) );
  BUF_X4 U98 ( .A(n19), .Z(n33) );
  BUF_X4 U99 ( .A(n13), .Z(n39) );
  BUF_X4 U100 ( .A(n9), .Z(n43) );
endmodule


module DECODE_UNIT_NB32_LS5 ( CLK, RST, FLUSH, DATAIN, IMM1, IMM2, BR_TYPE, 
        JMP, RI, US, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DEST_IN, HAZARD, 
        US_TO_EX, A, B, C, D, RT, RS, DEST_OUT );
  input [31:0] DATAIN;
  input [25:0] IMM1;
  input [31:0] IMM2;
  input [1:0] BR_TYPE;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [4:0] DEST_IN;
  output [31:0] A;
  output [31:0] B;
  output [31:0] C;
  output [31:0] D;
  output [4:0] RT;
  output [4:0] RS;
  output [4:0] DEST_OUT;
  input CLK, RST, FLUSH, JMP, RI, US, RD1, RD2, WR;
  output HAZARD, US_TO_EX;
  wire   n17, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n18, n19,
         n20, n21;
  wire   [31:0] OUT1;
  wire   [31:0] OUT2;
  wire   [31:0] EXT1;
  wire   [31:0] TO_IMM1;
  wire   [4:0] DEST_ADD;
  assign n17 = RST;

  register_file_NB32_RS32 reg_file ( .CLK(CLK), .RESET(n21), .RD1(RD1), .RD2(
        RD2), .WR(WR), .ADD_WR(ADD_WR), .ADD_RD1(ADD_RD1), .ADD_RD2(ADD_RD2), 
        .DATAIN(DATAIN), .HAZARD(HAZARD), .OUT1(OUT1), .OUT2(OUT2) );
  FD_INJ_NB32_4 reg_a ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(OUT1), .Q(
        A) );
  FD_INJ_NB32_3 reg_b ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(OUT2), .Q(
        B) );
  SIGN_EXT_NB32 exted ( .A(IMM1), .US(US), .JMP(JMP), .Y(EXT1) );
  FD_INJ_NB1_1 us_register ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(US), 
        .Q(US_TO_EX) );
  FD_INJ_NB32_2 imm_reg1 ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(TO_IMM1), .Q(C) );
  FD_INJ_NB32_1 imm_reg2 ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(IMM2), 
        .Q(D) );
  MUX21_generic_NB5 mux_dest ( .A(ADD_RD2), .B(DEST_IN), .SEL(RI), .Y(DEST_ADD) );
  FD_INJ_NB5_0 dest_reg ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(DEST_ADD), .Q(DEST_OUT) );
  FD_INJ_NB5_2 rs_reg ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(ADD_RD1), 
        .Q(RS) );
  FD_INJ_NB5_1 rt_reg ( .CK(CLK), .RESET(n21), .INJ_ZERO(FLUSH), .D(ADD_RD2), 
        .Q(RT) );
  NOR4_X1 U2 ( .A1(OUT1[23]), .A2(OUT1[22]), .A3(OUT1[21]), .A4(OUT1[20]), 
        .ZN(n9) );
  NOR4_X1 U3 ( .A1(OUT1[9]), .A2(OUT1[8]), .A3(OUT1[7]), .A4(OUT1[6]), .ZN(n13) );
  BUF_X2 U4 ( .A(n17), .Z(n21) );
  AND2_X1 U5 ( .A1(EXT1[25]), .A2(n19), .ZN(TO_IMM1[25]) );
  AND2_X1 U6 ( .A1(EXT1[26]), .A2(n19), .ZN(TO_IMM1[26]) );
  AND2_X1 U7 ( .A1(EXT1[27]), .A2(n19), .ZN(TO_IMM1[27]) );
  AND2_X1 U8 ( .A1(EXT1[28]), .A2(n18), .ZN(TO_IMM1[28]) );
  AND2_X1 U9 ( .A1(EXT1[29]), .A2(n18), .ZN(TO_IMM1[29]) );
  AND2_X1 U10 ( .A1(EXT1[30]), .A2(n18), .ZN(TO_IMM1[30]) );
  AND2_X1 U11 ( .A1(EXT1[31]), .A2(n18), .ZN(TO_IMM1[31]) );
  NOR4_X1 U12 ( .A1(OUT1[5]), .A2(OUT1[4]), .A3(OUT1[3]), .A4(OUT1[31]), .ZN(
        n12) );
  NOR4_X1 U13 ( .A1(OUT1[30]), .A2(OUT1[2]), .A3(OUT1[29]), .A4(OUT1[28]), 
        .ZN(n11) );
  NOR4_X1 U14 ( .A1(OUT1[27]), .A2(OUT1[26]), .A3(OUT1[25]), .A4(OUT1[24]), 
        .ZN(n10) );
  BUF_X1 U15 ( .A(n1), .Z(n19) );
  BUF_X1 U16 ( .A(n1), .Z(n18) );
  NAND4_X1 U17 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  NOR4_X1 U18 ( .A1(OUT1[12]), .A2(OUT1[11]), .A3(OUT1[10]), .A4(OUT1[0]), 
        .ZN(n6) );
  NOR4_X1 U19 ( .A1(OUT1[16]), .A2(OUT1[15]), .A3(OUT1[14]), .A4(OUT1[13]), 
        .ZN(n7) );
  NOR4_X1 U20 ( .A1(OUT1[1]), .A2(OUT1[19]), .A3(OUT1[18]), .A4(OUT1[17]), 
        .ZN(n8) );
  BUF_X1 U21 ( .A(n1), .Z(n20) );
  AND2_X1 U22 ( .A1(EXT1[0]), .A2(n20), .ZN(TO_IMM1[0]) );
  AND2_X1 U23 ( .A1(EXT1[1]), .A2(n19), .ZN(TO_IMM1[1]) );
  AND2_X1 U24 ( .A1(EXT1[2]), .A2(n18), .ZN(TO_IMM1[2]) );
  AND2_X1 U25 ( .A1(EXT1[10]), .A2(n20), .ZN(TO_IMM1[10]) );
  AND2_X1 U26 ( .A1(EXT1[11]), .A2(n20), .ZN(TO_IMM1[11]) );
  AND2_X1 U27 ( .A1(EXT1[12]), .A2(n20), .ZN(TO_IMM1[12]) );
  AND2_X1 U28 ( .A1(EXT1[13]), .A2(n20), .ZN(TO_IMM1[13]) );
  AND2_X1 U29 ( .A1(EXT1[14]), .A2(n20), .ZN(TO_IMM1[14]) );
  AND2_X1 U30 ( .A1(EXT1[15]), .A2(n20), .ZN(TO_IMM1[15]) );
  AND2_X1 U31 ( .A1(EXT1[16]), .A2(n20), .ZN(TO_IMM1[16]) );
  AND2_X1 U32 ( .A1(EXT1[17]), .A2(n19), .ZN(TO_IMM1[17]) );
  AND2_X1 U33 ( .A1(EXT1[18]), .A2(n19), .ZN(TO_IMM1[18]) );
  AND2_X1 U34 ( .A1(EXT1[19]), .A2(n19), .ZN(TO_IMM1[19]) );
  AND2_X1 U35 ( .A1(EXT1[20]), .A2(n19), .ZN(TO_IMM1[20]) );
  AND2_X1 U36 ( .A1(EXT1[21]), .A2(n19), .ZN(TO_IMM1[21]) );
  AND2_X1 U37 ( .A1(EXT1[22]), .A2(n19), .ZN(TO_IMM1[22]) );
  AND2_X1 U38 ( .A1(EXT1[23]), .A2(n19), .ZN(TO_IMM1[23]) );
  AND2_X1 U39 ( .A1(EXT1[24]), .A2(n19), .ZN(TO_IMM1[24]) );
  AND2_X1 U40 ( .A1(EXT1[9]), .A2(n18), .ZN(TO_IMM1[9]) );
  AND2_X1 U41 ( .A1(EXT1[3]), .A2(n18), .ZN(TO_IMM1[3]) );
  AND2_X1 U42 ( .A1(EXT1[4]), .A2(n18), .ZN(TO_IMM1[4]) );
  AND2_X1 U43 ( .A1(EXT1[5]), .A2(n18), .ZN(TO_IMM1[5]) );
  AND2_X1 U44 ( .A1(EXT1[6]), .A2(n18), .ZN(TO_IMM1[6]) );
  AND2_X1 U45 ( .A1(EXT1[7]), .A2(n18), .ZN(TO_IMM1[7]) );
  AND2_X1 U46 ( .A1(EXT1[8]), .A2(n18), .ZN(TO_IMM1[8]) );
  NAND2_X1 U47 ( .A1(n2), .A2(BR_TYPE[1]), .ZN(n1) );
  XNOR2_X1 U48 ( .A(BR_TYPE[0]), .B(n3), .ZN(n2) );
  NOR2_X1 U49 ( .A1(n4), .A2(n5), .ZN(n3) );
  NAND4_X1 U50 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(n4) );
endmodule


module FETCH_UNIT_NB32_LS5 ( CLK, STALL, RST, RST_DEC, PC_SEL, JB_INST, 
        IRAM_OUT, FUNC, OPCODE, CURR_PC, NPC, INST_OUT, MISS_HIT );
  input [31:0] JB_INST;
  input [31:0] IRAM_OUT;
  output [10:0] FUNC;
  output [5:0] OPCODE;
  output [31:0] CURR_PC;
  output [31:0] NPC;
  output [31:0] INST_OUT;
  output [1:0] MISS_HIT;
  input CLK, STALL, RST, RST_DEC, PC_SEL;
  wire   \IRAM_OUT[10] , \IRAM_OUT[9] , \IRAM_OUT[8] , \IRAM_OUT[7] ,
         \IRAM_OUT[6] , \IRAM_OUT[5] , \IRAM_OUT[4] , \IRAM_OUT[3] ,
         \IRAM_OUT[2] , \IRAM_OUT[1] , \IRAM_OUT[0] , \IRAM_OUT[31] ,
         \IRAM_OUT[30] , \IRAM_OUT[29] , \IRAM_OUT[28] , \IRAM_OUT[27] ,
         \IRAM_OUT[26] , TMP_RST, n7, n8, n9;
  wire   [31:0] NEXT_PC;
  wire   [31:0] NEW_PC;
  wire   [31:0] TMP_INST_OUT;
  wire   [31:0] PRED;
  assign FUNC[10] = \IRAM_OUT[10] ;
  assign \IRAM_OUT[10]  = IRAM_OUT[10];
  assign FUNC[9] = \IRAM_OUT[9] ;
  assign \IRAM_OUT[9]  = IRAM_OUT[9];
  assign FUNC[8] = \IRAM_OUT[8] ;
  assign \IRAM_OUT[8]  = IRAM_OUT[8];
  assign FUNC[7] = \IRAM_OUT[7] ;
  assign \IRAM_OUT[7]  = IRAM_OUT[7];
  assign FUNC[6] = \IRAM_OUT[6] ;
  assign \IRAM_OUT[6]  = IRAM_OUT[6];
  assign FUNC[5] = \IRAM_OUT[5] ;
  assign \IRAM_OUT[5]  = IRAM_OUT[5];
  assign FUNC[4] = \IRAM_OUT[4] ;
  assign \IRAM_OUT[4]  = IRAM_OUT[4];
  assign FUNC[3] = \IRAM_OUT[3] ;
  assign \IRAM_OUT[3]  = IRAM_OUT[3];
  assign FUNC[2] = \IRAM_OUT[2] ;
  assign \IRAM_OUT[2]  = IRAM_OUT[2];
  assign FUNC[1] = \IRAM_OUT[1] ;
  assign \IRAM_OUT[1]  = IRAM_OUT[1];
  assign FUNC[0] = \IRAM_OUT[0] ;
  assign \IRAM_OUT[0]  = IRAM_OUT[0];
  assign OPCODE[5] = \IRAM_OUT[31] ;
  assign \IRAM_OUT[31]  = IRAM_OUT[31];
  assign OPCODE[4] = \IRAM_OUT[30] ;
  assign \IRAM_OUT[30]  = IRAM_OUT[30];
  assign OPCODE[3] = \IRAM_OUT[29] ;
  assign \IRAM_OUT[29]  = IRAM_OUT[29];
  assign OPCODE[2] = \IRAM_OUT[28] ;
  assign \IRAM_OUT[28]  = IRAM_OUT[28];
  assign OPCODE[1] = \IRAM_OUT[27] ;
  assign \IRAM_OUT[27]  = IRAM_OUT[27];
  assign OPCODE[0] = \IRAM_OUT[26] ;
  assign \IRAM_OUT[26]  = IRAM_OUT[26];

  DFF_X1 TMP_RST_reg ( .D(RST), .CK(CLK), .Q(TMP_RST) );
  FD_INJ_NB32_0 N_PC ( .CK(CLK), .RESET(RST), .INJ_ZERO(n9), .D(NEXT_PC), .Q(
        NPC) );
  BP_NB32_BP_LEN4 BP_UNIT ( .CLK(CLK), .RST(RST), .EX_PC(JB_INST), .CURR_PC(
        CURR_PC), .NEXT_PC(NEXT_PC), .NEW_PC(NEW_PC), .INST(TMP_INST_OUT), 
        .MISS_HIT(MISS_HIT), .PRED(PRED) );
  FD_NB32_0 PC ( .CK(CLK), .RESET(TMP_RST), .D(PRED), .Q(CURR_PC) );
  MUX21_generic_NB32_0 flush_mux ( .A({\IRAM_OUT[31] , \IRAM_OUT[30] , 
        \IRAM_OUT[29] , \IRAM_OUT[28] , \IRAM_OUT[27] , \IRAM_OUT[26] , 
        IRAM_OUT[25:11], \IRAM_OUT[10] , \IRAM_OUT[9] , \IRAM_OUT[8] , 
        \IRAM_OUT[7] , \IRAM_OUT[6] , \IRAM_OUT[5] , \IRAM_OUT[4] , 
        \IRAM_OUT[3] , \IRAM_OUT[2] , \IRAM_OUT[1] , \IRAM_OUT[0] }), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n7), .Y(TMP_INST_OUT)
         );
  FD_NB32_5 INST ( .CK(CLK), .RESET(RST), .D(TMP_INST_OUT), .Q(INST_OUT) );
  MUX21_generic_NB32_4 pc_mux ( .A(JB_INST), .B(NEXT_PC), .SEL(PC_SEL), .Y(
        NEW_PC) );
  FETCH_UNIT_NB32_LS5_DW01_add_0 add_123 ( .A(CURR_PC), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NEXT_PC) );
  CLKBUF_X1 U5 ( .A(n7), .Z(n9) );
  AOI21_X1 U7 ( .B1(MISS_HIT[0]), .B2(MISS_HIT[1]), .A(n8), .ZN(n7) );
  INV_X1 U8 ( .A(STALL), .ZN(n8) );
endmodule


module DLX_CU ( CLK, RST, OPCODE, FUNC, FLUSH, STALL, JMP, RI, BR_TYPE, RD1, 
        RD2, US, MUX1_SEL, MUX2_SEL, UN_SEL, OP_SEL, PC_SEL, RW, D_TYPE, WR, 
        MEM_ALU_SEL, INST_T_EX, .INST_EX({\INST_EX[1] , \INST_EX[0] }), 
    .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }) );
  input [5:0] OPCODE;
  input [10:0] FUNC;
  output [1:0] BR_TYPE;
  output [2:0] UN_SEL;
  output [3:0] OP_SEL;
  output [1:0] D_TYPE;
  input CLK, RST, FLUSH;
  output STALL, JMP, RI, RD1, RD2, US, MUX1_SEL, MUX2_SEL, PC_SEL, RW, WR,
         MEM_ALU_SEL, INST_T_EX, \INST_EX[1] , \INST_EX[0] , \INST_MEM[1] ,
         \INST_MEM[0] ;
  wire   \TMP1E[0] , \TMP2E[0] , \TMP5E[0] , \TMP11M[0] , \TMP12M[0] ,
         \TMP11W[0] , \TMP21W[0] , \TMP12W[0] , \TMP22W[0] , \TMP13W[0] ,
         \TMP23W[0] , \INST_TMP[0] , \INST_TMP1[0] , n8, n179, n182, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n180, n181, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n207, n208,
         n209, n206, n210;
  wire   [5:0] OPCODE1;
  wire   [5:0] OPCODE2;
  wire   [5:0] OPCODE3;
  wire   [10:0] FUNC1;
  wire   [1:0] INST;
  wire   [1:0] NEXT_INST;
  wire   [21:0] cw;
  wire   [2:0] TMP3E;
  wire   [3:0] TMP4E;
  wire   [1:0] TMP21M;
  wire   [1:0] TMP22M;
  wire   [1:0] INST1;
  assign n182 = RST;

  DFFR_X1 \INST_reg[1]  ( .D(NEXT_INST[1]), .CK(CLK), .RN(n210), .Q(INST[1]), 
        .QN(n8) );
  DFFR_X1 \INST1_reg[1]  ( .D(INST[1]), .CK(CLK), .RN(n210), .Q(INST1[1]) );
  DFFR_X1 \INST1_reg[0]  ( .D(INST[0]), .CK(CLK), .RN(n210), .Q(INST1[0]) );
  DFFR_X1 \INST2_reg[1]  ( .D(INST1[1]), .CK(CLK), .RN(n210), .Q(INST_EX[1])
         );
  DFFR_X1 \INST2_reg[0]  ( .D(INST1[0]), .CK(CLK), .RN(n210), .Q(INST_EX[0])
         );
  DFFR_X1 \INST3_reg[1]  ( .D(INST_EX[1]), .CK(CLK), .RN(n210), .Q(INST_MEM[1]) );
  DFFR_X1 \INST3_reg[0]  ( .D(INST_EX[0]), .CK(CLK), .RN(n210), .Q(INST_MEM[0]) );
  DFFR_X1 \INST_reg[0]  ( .D(NEXT_INST[0]), .CK(CLK), .RN(n210), .Q(INST[0]), 
        .QN(n179) );
  NAND3_X1 U166 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n62) );
  NAND3_X1 U167 ( .A1(n136), .A2(n137), .A3(n138), .ZN(n135) );
  NAND3_X1 U168 ( .A1(n111), .A2(n103), .A3(n118), .ZN(STALL) );
  NAND3_X1 U169 ( .A1(n158), .A2(n148), .A3(n165), .ZN(n164) );
  NAND3_X1 U170 ( .A1(n167), .A2(n168), .A3(n169), .ZN(n134) );
  NAND3_X1 U171 ( .A1(FUNC[2]), .A2(n173), .A3(n170), .ZN(n67) );
  NAND3_X1 U172 ( .A1(n173), .A2(n167), .A3(n100), .ZN(n70) );
  NAND3_X1 U173 ( .A1(n173), .A2(n167), .A3(n132), .ZN(n77) );
  NAND3_X1 U174 ( .A1(FUNC[3]), .A2(n167), .A3(n169), .ZN(n65) );
  NAND3_X1 U175 ( .A1(FUNC[2]), .A2(n173), .A3(n133), .ZN(n81) );
  NAND3_X1 U176 ( .A1(n184), .A2(n185), .A3(n86), .ZN(n183) );
  NAND3_X1 U177 ( .A1(n86), .A2(n185), .A3(n186), .ZN(n116) );
  NAND3_X1 U178 ( .A1(n119), .A2(n115), .A3(n113), .ZN(n104) );
  NAND3_X1 U179 ( .A1(n108), .A2(OPCODE[5]), .A3(n191), .ZN(n115) );
  NAND3_X1 U180 ( .A1(OPCODE[1]), .A2(n195), .A3(n185), .ZN(n154) );
  NAND3_X1 U181 ( .A1(n190), .A2(OPCODE[3]), .A3(OPCODE[1]), .ZN(n93) );
  NAND3_X1 U182 ( .A1(n185), .A2(n195), .A3(n53), .ZN(n128) );
  NAND3_X1 U183 ( .A1(OPCODE[3]), .A2(n201), .A3(n185), .ZN(n84) );
  NAND3_X1 U184 ( .A1(OPCODE1[1]), .A2(n208), .A3(n209), .ZN(n205) );
  NAND3_X1 U185 ( .A1(n83), .A2(n200), .A3(n184), .ZN(n180) );
  FD_NB6_0 OPPP1 ( .CK(CLK), .RESET(n206), .D(OPCODE), .Q(OPCODE1) );
  FD_NB6_3 OPPP2 ( .CK(CLK), .RESET(n206), .D(OPCODE1), .Q(OPCODE2) );
  FD_NB6_2 OPPP3 ( .CK(CLK), .RESET(n206), .D(OPCODE2), .Q(OPCODE3) );
  FD_NB6_1 OPPP4 ( .CK(CLK), .RESET(n206), .D(OPCODE3) );
  FD_NB11_0 FUNPP1 ( .CK(CLK), .RESET(n206), .D(FUNC), .Q(FUNC1) );
  FD_NB11_1 FUNPP2 ( .CK(CLK), .RESET(n206), .D(FUNC1) );
  FD_NB1_0 pipe1_JMP ( .CK(CLK), .RESET(n210), .D(cw[21]), .Q(JMP) );
  FD_NB1_22 pipe1_RI ( .CK(CLK), .RESET(n210), .D(cw[20]), .Q(RI) );
  FD_NB2_0 pipe1_BR ( .CK(CLK), .RESET(n210), .D(cw[19:18]), .Q(BR_TYPE) );
  FD_NB1_21 pipe1_RD1 ( .CK(CLK), .RESET(n210), .D(cw[17]), .Q(RD1) );
  FD_NB1_20 pipe1_RD2 ( .CK(CLK), .RESET(n210), .D(cw[16]), .Q(RD2) );
  FD_NB1_19 pipe1_US ( .CK(CLK), .RESET(n210), .D(cw[15]), .Q(US) );
  FD_NB1_18 pipe1_MX1 ( .CK(CLK), .RESET(n210), .D(cw[14]), .Q(\TMP1E[0] ) );
  FD_NB1_17 pipe1_MX2 ( .CK(CLK), .RESET(n210), .D(cw[13]), .Q(\TMP2E[0] ) );
  FD_NB3_0 pipe1_UN ( .CK(CLK), .RESET(n210), .D(cw[12:10]), .Q(TMP3E) );
  FD_NB4_0 pipe1_OP ( .CK(CLK), .RESET(n206), .D(cw[9:6]), .Q(TMP4E) );
  FD_NB1_16 pipe1_PC ( .CK(CLK), .RESET(n210), .D(cw[5]), .Q(\TMP5E[0] ) );
  FD_NB1_15 pipe2_MX1 ( .CK(CLK), .RESET(n210), .D(\TMP1E[0] ), .Q(MUX1_SEL)
         );
  FD_NB1_14 pipe2_MX2 ( .CK(CLK), .RESET(n210), .D(\TMP2E[0] ), .Q(MUX2_SEL)
         );
  FD_NB3_1 pipe2_UN ( .CK(CLK), .RESET(n210), .D(TMP3E), .Q(UN_SEL) );
  FD_NB4_1 pipe2_OP ( .CK(CLK), .RESET(n206), .D(TMP4E), .Q(OP_SEL) );
  FD_NB1_13 pipe2_PC ( .CK(CLK), .RESET(n210), .D(\TMP5E[0] ), .Q(PC_SEL) );
  FD_NB1_12 pipe1_RW ( .CK(CLK), .RESET(n210), .D(cw[4]), .Q(\TMP11M[0] ) );
  FD_NB2_3 pipe1_DT ( .CK(CLK), .RESET(n210), .D(cw[3:2]), .Q(TMP21M) );
  FD_NB1_11 pipe2_RW ( .CK(CLK), .RESET(n210), .D(\TMP11M[0] ), .Q(\TMP12M[0] ) );
  FD_NB2_2 pipe2_DT ( .CK(CLK), .RESET(n210), .D(TMP21M), .Q(TMP22M) );
  FD_NB1_10 pipe3_RW ( .CK(CLK), .RESET(n210), .D(\TMP12M[0] ), .Q(RW) );
  FD_NB2_1 pipe3_DT ( .CK(CLK), .RESET(n210), .D(TMP22M), .Q(D_TYPE) );
  FD_INJ_NB1_0 pipe1_WR ( .CK(CLK), .RESET(n210), .INJ_ZERO(FLUSH), .D(cw[1]), 
        .Q(\TMP11W[0] ) );
  FD_NB1_9 pipe1_MM ( .CK(CLK), .RESET(n210), .D(cw[0]), .Q(\TMP21W[0] ) );
  FD_INJ_NB1_2 pipe2_WR ( .CK(CLK), .RESET(FLUSH), .INJ_ZERO(n210), .D(
        \TMP11W[0] ), .Q(\TMP12W[0] ) );
  FD_NB1_8 pipe2_MM ( .CK(CLK), .RESET(n210), .D(\TMP21W[0] ), .Q(\TMP22W[0] )
         );
  FD_NB1_7 pipe3_WR ( .CK(CLK), .RESET(n210), .D(\TMP12W[0] ), .Q(\TMP13W[0] )
         );
  FD_NB1_6 pipe3_MM ( .CK(CLK), .RESET(n210), .D(\TMP22W[0] ), .Q(\TMP23W[0] )
         );
  FD_NB1_5 pipe4_WR ( .CK(CLK), .RESET(n210), .D(\TMP13W[0] ), .Q(WR) );
  FD_NB1_4 pipe4_MM ( .CK(CLK), .RESET(n210), .D(\TMP23W[0] ), .Q(MEM_ALU_SEL)
         );
  FD_NB1_3 pipe1_INST ( .CK(CLK), .RESET(n210), .D(\INST_TMP[0] ), .Q(
        \INST_TMP1[0] ) );
  FD_NB1_2 pipe2_INST ( .CK(CLK), .RESET(n210), .D(\INST_TMP1[0] ), .Q(
        INST_T_EX) );
  NOR4_X1 U3 ( .A1(n167), .A2(FUNC[3]), .A3(FUNC[4]), .A4(FUNC[5]), .ZN(n101)
         );
  NOR4_X1 U4 ( .A1(FUNC[6]), .A2(FUNC[10]), .A3(n180), .A4(n181), .ZN(n75) );
  INV_X1 U5 ( .A(n111), .ZN(cw[20]) );
  INV_X1 U6 ( .A(n103), .ZN(cw[5]) );
  NAND2_X1 U7 ( .A1(n86), .A2(n140), .ZN(n111) );
  NOR2_X1 U8 ( .A1(n102), .A2(n171), .ZN(n158) );
  INV_X1 U9 ( .A(n130), .ZN(n171) );
  NOR2_X1 U10 ( .A1(cw[19]), .A2(cw[21]), .ZN(n103) );
  INV_X1 U11 ( .A(n128), .ZN(n151) );
  NAND2_X1 U12 ( .A1(n162), .A2(n86), .ZN(n118) );
  INV_X1 U13 ( .A(n137), .ZN(n162) );
  AOI21_X1 U14 ( .B1(n89), .B2(n73), .A(n90), .ZN(n72) );
  NAND2_X1 U15 ( .A1(n139), .A2(n73), .ZN(n136) );
  INV_X1 U16 ( .A(n134), .ZN(n99) );
  INV_X1 U17 ( .A(n163), .ZN(n139) );
  INV_X1 U18 ( .A(cw[21]), .ZN(n142) );
  INV_X1 U19 ( .A(n180), .ZN(\INST_TMP[0] ) );
  INV_X1 U20 ( .A(n116), .ZN(cw[18]) );
  NAND2_X1 U21 ( .A1(n117), .A2(n118), .ZN(cw[16]) );
  INV_X1 U22 ( .A(cw[4]), .ZN(n117) );
  OR2_X1 U23 ( .A1(cw[14]), .A2(cw[19]), .ZN(cw[17]) );
  AND2_X1 U24 ( .A1(n104), .A2(n86), .ZN(cw[3]) );
  NAND4_X1 U25 ( .A1(n110), .A2(n125), .A3(n187), .A4(n188), .ZN(n140) );
  AND3_X1 U26 ( .A1(n147), .A2(n60), .A3(n59), .ZN(n187) );
  NOR4_X1 U27 ( .A1(n151), .A2(n96), .A3(n189), .A4(n104), .ZN(n188) );
  INV_X1 U28 ( .A(n114), .ZN(n189) );
  OAI221_X1 U29 ( .B1(n194), .B2(n84), .C1(n92), .C2(n196), .A(n197), .ZN(n56)
         );
  INV_X1 U30 ( .A(n123), .ZN(n197) );
  NOR2_X1 U31 ( .A1(n53), .A2(n73), .ZN(n194) );
  INV_X1 U32 ( .A(n196), .ZN(n73) );
  INV_X1 U33 ( .A(n93), .ZN(n107) );
  OR2_X1 U34 ( .A1(n157), .A2(n54), .ZN(n96) );
  OR2_X1 U35 ( .A1(n56), .A2(n193), .ZN(n157) );
  AOI21_X1 U36 ( .B1(n154), .B2(n125), .A(n194), .ZN(n193) );
  OR2_X1 U37 ( .A1(cw[0]), .A2(n112), .ZN(cw[1]) );
  AOI21_X1 U38 ( .B1(n113), .B2(n106), .A(n52), .ZN(n112) );
  OAI21_X1 U39 ( .B1(n170), .B2(n100), .A(n101), .ZN(n130) );
  INV_X1 U40 ( .A(n52), .ZN(n86) );
  NOR2_X1 U41 ( .A1(n163), .A2(n52), .ZN(cw[21]) );
  AOI21_X1 U42 ( .B1(n190), .B2(n184), .A(n122), .ZN(n114) );
  AOI21_X1 U43 ( .B1(n190), .B2(n186), .A(n124), .ZN(n113) );
  NAND4_X1 U44 ( .A1(n81), .A2(n76), .A3(n87), .A4(n172), .ZN(n102) );
  AND4_X1 U45 ( .A1(n65), .A2(n153), .A3(n68), .A4(n67), .ZN(n172) );
  NAND2_X1 U46 ( .A1(n75), .A2(n164), .ZN(n137) );
  AND3_X1 U47 ( .A1(n66), .A2(n134), .A3(n69), .ZN(n165) );
  NAND2_X1 U48 ( .A1(n101), .A2(n132), .ZN(n153) );
  OAI21_X1 U49 ( .B1(n192), .B2(n107), .A(n108), .ZN(n119) );
  NAND2_X1 U50 ( .A1(n191), .A2(n200), .ZN(n163) );
  INV_X1 U51 ( .A(n91), .ZN(n125) );
  OR2_X1 U52 ( .A1(n203), .A2(n84), .ZN(n60) );
  OR2_X1 U53 ( .A1(n126), .A2(n84), .ZN(n59) );
  INV_X1 U54 ( .A(n64), .ZN(n100) );
  INV_X1 U55 ( .A(n54), .ZN(n92) );
  NAND2_X1 U56 ( .A1(n192), .A2(n204), .ZN(n110) );
  NAND2_X1 U57 ( .A1(n170), .A2(n166), .ZN(n66) );
  NAND2_X1 U58 ( .A1(n116), .A2(n183), .ZN(cw[19]) );
  NAND2_X1 U59 ( .A1(n166), .A2(n133), .ZN(n69) );
  INV_X1 U60 ( .A(n126), .ZN(n108) );
  NAND2_X1 U61 ( .A1(n174), .A2(n170), .ZN(n68) );
  NAND2_X1 U62 ( .A1(n64), .A2(n80), .ZN(n98) );
  INV_X1 U63 ( .A(n80), .ZN(n132) );
  NAND2_X1 U64 ( .A1(n174), .A2(n133), .ZN(n76) );
  INV_X1 U65 ( .A(n199), .ZN(n82) );
  INV_X1 U66 ( .A(n175), .ZN(n87) );
  OAI211_X1 U67 ( .C1(n176), .C2(n65), .A(n77), .B(n70), .ZN(n175) );
  NOR2_X1 U68 ( .A1(n133), .A2(n98), .ZN(n176) );
  NAND2_X1 U69 ( .A1(n166), .A2(n100), .ZN(n148) );
  INV_X1 U70 ( .A(n204), .ZN(n203) );
  NOR2_X1 U71 ( .A1(n149), .A2(n52), .ZN(cw[11]) );
  AOI211_X1 U72 ( .C1(n150), .C2(n73), .A(n151), .B(n152), .ZN(n149) );
  INV_X1 U73 ( .A(n154), .ZN(n150) );
  AOI21_X1 U74 ( .B1(n130), .B2(n153), .A(n58), .ZN(n152) );
  OAI221_X1 U75 ( .B1(n52), .B2(n136), .C1(n141), .C2(n142), .A(n118), .ZN(
        cw[13]) );
  INV_X1 U76 ( .A(n53), .ZN(n141) );
  OAI21_X1 U77 ( .B1(n126), .B2(n163), .A(n136), .ZN(n145) );
  INV_X1 U78 ( .A(n75), .ZN(n58) );
  OAI211_X1 U79 ( .C1(n146), .C2(n58), .A(n147), .B(n59), .ZN(n90) );
  AND2_X1 U80 ( .A1(n148), .A2(n69), .ZN(n146) );
  NOR2_X1 U81 ( .A1(n143), .A2(n52), .ZN(cw[12]) );
  NOR3_X1 U82 ( .A1(n144), .A2(n90), .A3(n145), .ZN(n143) );
  OAI21_X1 U83 ( .B1(n58), .B2(n66), .A(n60), .ZN(n144) );
  NOR2_X1 U84 ( .A1(n155), .A2(n52), .ZN(cw[10]) );
  NOR3_X1 U85 ( .A1(n156), .A2(n157), .A3(n145), .ZN(n155) );
  OAI21_X1 U86 ( .B1(n158), .B2(n58), .A(n128), .ZN(n156) );
  AOI21_X1 U87 ( .B1(n110), .B2(n119), .A(n52), .ZN(cw[4]) );
  NOR2_X1 U88 ( .A1(n51), .A2(n52), .ZN(cw[9]) );
  AOI211_X1 U89 ( .C1(n53), .C2(n54), .A(n55), .B(n56), .ZN(n51) );
  OAI211_X1 U90 ( .C1(n57), .C2(n58), .A(n59), .B(n60), .ZN(n55) );
  NOR3_X1 U91 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n57) );
  OAI21_X1 U92 ( .B1(n64), .B2(n65), .A(n66), .ZN(n63) );
  NAND4_X1 U93 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(n61) );
  AOI21_X1 U94 ( .B1(n105), .B2(n106), .A(n52), .ZN(cw[2]) );
  AOI21_X1 U95 ( .B1(n107), .B2(n108), .A(n109), .ZN(n105) );
  INV_X1 U96 ( .A(n110), .ZN(n109) );
  AOI21_X1 U97 ( .B1(n71), .B2(n72), .A(n52), .ZN(cw[8]) );
  AOI22_X1 U98 ( .A1(n73), .A2(n74), .B1(n75), .B2(n62), .ZN(n71) );
  OAI21_X1 U99 ( .B1(n82), .B2(n83), .A(n84), .ZN(n74) );
  NAND2_X1 U100 ( .A1(n92), .A2(n93), .ZN(n89) );
  OAI21_X1 U101 ( .B1(n205), .B2(INST[0]), .A(n142), .ZN(NEXT_INST[1]) );
  NOR2_X1 U102 ( .A1(n120), .A2(n52), .ZN(cw[15]) );
  NOR4_X1 U103 ( .A1(n121), .A2(n122), .A3(n123), .A4(n124), .ZN(n120) );
  OAI221_X1 U104 ( .B1(n125), .B2(n126), .C1(n127), .C2(n58), .A(n128), .ZN(
        n121) );
  AND4_X1 U105 ( .A1(n129), .A2(n67), .A3(n130), .A4(n70), .ZN(n127) );
  NOR2_X1 U106 ( .A1(n94), .A2(n52), .ZN(cw[6]) );
  AOI21_X1 U107 ( .B1(n75), .B2(n95), .A(n96), .ZN(n94) );
  INV_X1 U108 ( .A(n97), .ZN(n95) );
  AOI221_X1 U109 ( .B1(n98), .B2(n99), .C1(n100), .C2(n101), .A(n102), .ZN(n97) );
  AND2_X1 U110 ( .A1(n114), .A2(n115), .ZN(n106) );
  AND3_X1 U111 ( .A1(n81), .A2(n77), .A3(n131), .ZN(n129) );
  OAI21_X1 U112 ( .B1(n132), .B2(n133), .A(n99), .ZN(n131) );
  AND2_X1 U113 ( .A1(n86), .A2(n135), .ZN(cw[14]) );
  AOI21_X1 U114 ( .B1(n139), .B2(n53), .A(n140), .ZN(n138) );
  INV_X1 U115 ( .A(n159), .ZN(cw[0]) );
  OAI21_X1 U116 ( .B1(n160), .B2(n161), .A(n86), .ZN(n159) );
  NAND4_X1 U117 ( .A1(n125), .A2(n147), .A3(n59), .A4(n60), .ZN(n160) );
  OR4_X1 U118 ( .A1(n145), .A2(n96), .A3(n162), .A4(n151), .ZN(n161) );
  INV_X1 U119 ( .A(n79), .ZN(n78) );
  OAI21_X1 U120 ( .B1(n65), .B2(n80), .A(n81), .ZN(n79) );
  AND2_X1 U121 ( .A1(n85), .A2(n86), .ZN(cw[7]) );
  OAI211_X1 U122 ( .C1(n58), .C2(n87), .A(n88), .B(n72), .ZN(n85) );
  AOI22_X1 U123 ( .A1(n91), .A2(n73), .B1(n89), .B2(n53), .ZN(n88) );
  NOR2_X1 U124 ( .A1(n202), .A2(OPCODE[0]), .ZN(n53) );
  NOR3_X1 U125 ( .A1(n195), .A2(OPCODE[1]), .A3(n200), .ZN(n199) );
  NOR2_X1 U126 ( .A1(n200), .A2(OPCODE[2]), .ZN(n190) );
  NOR2_X1 U127 ( .A1(n198), .A2(n194), .ZN(n123) );
  AOI21_X1 U128 ( .B1(n199), .B2(OPCODE[2]), .A(n107), .ZN(n198) );
  INV_X1 U129 ( .A(OPCODE[3]), .ZN(n195) );
  INV_X1 U130 ( .A(OPCODE[5]), .ZN(n200) );
  NAND2_X1 U131 ( .A1(OPCODE[4]), .A2(OPCODE[0]), .ZN(n196) );
  INV_X1 U132 ( .A(OPCODE[4]), .ZN(n202) );
  OR3_X1 U133 ( .A1(FUNC[9]), .A2(FUNC[8]), .A3(FUNC[7]), .ZN(n181) );
  NOR4_X1 U134 ( .A1(n201), .A2(n195), .A3(OPCODE[2]), .A4(OPCODE[5]), .ZN(n54) );
  NAND2_X1 U135 ( .A1(n8), .A2(INST[0]), .ZN(n52) );
  NOR3_X1 U136 ( .A1(OPCODE[1]), .A2(OPCODE[3]), .A3(n203), .ZN(n184) );
  NOR2_X1 U137 ( .A1(n177), .A2(FUNC[1]), .ZN(n133) );
  NOR3_X1 U138 ( .A1(OPCODE[1]), .A2(OPCODE[3]), .A3(n126), .ZN(n186) );
  NOR3_X1 U139 ( .A1(OPCODE[2]), .A2(OPCODE[5]), .A3(n195), .ZN(n91) );
  NOR2_X1 U140 ( .A1(n83), .A2(OPCODE[5]), .ZN(n185) );
  NOR2_X1 U141 ( .A1(FUNC[1]), .A2(FUNC[0]), .ZN(n170) );
  NOR3_X1 U142 ( .A1(OPCODE[2]), .A2(OPCODE[3]), .A3(n201), .ZN(n191) );
  NOR2_X1 U143 ( .A1(OPCODE[4]), .A2(OPCODE[0]), .ZN(n204) );
  NAND4_X1 U144 ( .A1(n204), .A2(n185), .A3(OPCODE[1]), .A4(OPCODE[3]), .ZN(
        n147) );
  NOR2_X1 U145 ( .A1(n178), .A2(FUNC[4]), .ZN(n169) );
  INV_X1 U146 ( .A(FUNC[5]), .ZN(n178) );
  NAND2_X1 U147 ( .A1(OPCODE[0]), .A2(n202), .ZN(n126) );
  NOR2_X1 U148 ( .A1(n82), .A2(OPCODE[2]), .ZN(n192) );
  NAND2_X1 U149 ( .A1(FUNC[0]), .A2(FUNC[1]), .ZN(n80) );
  AND3_X1 U150 ( .A1(n169), .A2(n168), .A3(FUNC[2]), .ZN(n166) );
  NAND2_X1 U151 ( .A1(FUNC[1]), .A2(n177), .ZN(n64) );
  INV_X1 U152 ( .A(FUNC[2]), .ZN(n167) );
  AND3_X1 U153 ( .A1(FUNC[4]), .A2(FUNC[3]), .A3(FUNC[5]), .ZN(n173) );
  AND3_X1 U154 ( .A1(OPCODE[2]), .A2(OPCODE[5]), .A3(n186), .ZN(n124) );
  AND3_X1 U155 ( .A1(OPCODE[2]), .A2(OPCODE[5]), .A3(n184), .ZN(n122) );
  AND3_X1 U156 ( .A1(n169), .A2(FUNC[3]), .A3(FUNC[2]), .ZN(n174) );
  INV_X1 U157 ( .A(OPCODE[1]), .ZN(n201) );
  INV_X1 U158 ( .A(OPCODE[2]), .ZN(n83) );
  INV_X1 U159 ( .A(FUNC[0]), .ZN(n177) );
  INV_X1 U160 ( .A(FUNC[3]), .ZN(n168) );
  BUF_X2 U161 ( .A(n182), .Z(n210) );
  INV_X1 U162 ( .A(OPCODE1[2]), .ZN(n208) );
  NOR3_X1 U163 ( .A1(OPCODE1[3]), .A2(n8), .A3(OPCODE1[5]), .ZN(n209) );
  INV_X1 U164 ( .A(n207), .ZN(NEXT_INST[0]) );
  AOI22_X1 U165 ( .A1(n163), .A2(n8), .B1(n205), .B2(n179), .ZN(n207) );
  CLKBUF_X3 U186 ( .A(n182), .Z(n206) );
endmodule


module DATAPATH_NB32_LS5_OPC6_FN11 ( CLK, STALL, RST, .INST_EX({\INST_EX[1] , 
        \INST_EX[0] }), .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }), INST_T_EX, 
        JMP, RI, RD1, RD2, WR, PC_SEL, MEM_ALU_SEL, US, MUX1_SEL, MUX2_SEL, 
        BR_TYPE, UN_SEL, OP_SEL, IRAM_OUT, EXT_MEM_IN, FLUSH, US_MEM, HAZARD, 
        EXT_MEM_ADD, EXT_MEM_DATA, CURR_PC, FUNC, OP_CODE );
  input [1:0] BR_TYPE;
  input [2:0] UN_SEL;
  input [3:0] OP_SEL;
  input [31:0] IRAM_OUT;
  input [31:0] EXT_MEM_IN;
  output [4:0] EXT_MEM_ADD;
  output [31:0] EXT_MEM_DATA;
  output [31:0] CURR_PC;
  output [10:0] FUNC;
  output [5:0] OP_CODE;
  input CLK, STALL, RST, \INST_EX[1] , \INST_EX[0] , \INST_MEM[1] ,
         \INST_MEM[0] , INST_T_EX, JMP, RI, RD1, RD2, WR, PC_SEL, MEM_ALU_SEL,
         US, MUX1_SEL, MUX2_SEL;
  output FLUSH, US_MEM, HAZARD;
  wire   US_TO_EX, n6, n5;
  wire   [1:0] MISS_HIT;
  wire   [31:0] TEMP_PC;
  wire   [31:0] NPC;
  wire   [25:0] INST;
  wire   [31:0] DATA_WB;
  wire   [4:0] DEST_FROM_WRBU;
  wire   [31:0] A;
  wire   [31:0] B;
  wire   [31:0] C;
  wire   [31:0] D;
  wire   [4:0] RT;
  wire   [4:0] RS;
  wire   [4:0] DEST_FROM_DECU;
  wire   [1:0] FW_MUX1_SEL;
  wire   [1:0] FW_MUX2_SEL;
  wire   [31:5] ALU_OUT;
  wire   [4:0] DEST_FROM_EXEU;
  wire   [31:0] ALU_TO_WB;
  wire   [31:0] TMP_MEM;
  wire   [4:0] DEST_FROM_MEMU;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5;

  FETCH_UNIT_NB32_LS5 ife_unit ( .CLK(CLK), .STALL(STALL), .RST(RST), 
        .RST_DEC(RST), .PC_SEL(PC_SEL), .JB_INST(TEMP_PC), .IRAM_OUT(IRAM_OUT), 
        .FUNC(FUNC), .OPCODE(OP_CODE), .CURR_PC(CURR_PC), .NPC(NPC), 
        .INST_OUT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, INST}), .MISS_HIT(
        MISS_HIT) );
  DECODE_UNIT_NB32_LS5 dec_unit ( .CLK(CLK), .RST(RST), .FLUSH(FLUSH), 
        .DATAIN(DATA_WB), .IMM1(INST), .IMM2(NPC), .BR_TYPE(BR_TYPE), .JMP(JMP), .RI(RI), .US(US), .RD1(RD1), .RD2(RD2), .WR(WR), .ADD_WR(DEST_FROM_WRBU), 
        .ADD_RD1(INST[25:21]), .ADD_RD2(INST[20:16]), .DEST_IN(INST[15:11]), 
        .HAZARD(HAZARD), .US_TO_EX(US_TO_EX), .A(A), .B(B), .C(C), .D(D), .RT(
        RT), .RS(RS), .DEST_OUT(DEST_FROM_DECU) );
  EXECUTION_UNIT_NB32_LS5 exe_unit ( .FW_MUX1_SEL(FW_MUX1_SEL), .FW_MUX2_SEL(
        FW_MUX2_SEL), .FW_EX({ALU_OUT, EXT_MEM_ADD}), .FW_MEM(DATA_WB), .A(A), 
        .B(B), .C(C), .D(D), .DEST_IN(DEST_FROM_DECU), .CLK(CLK), .RST(RST), 
        .US(US_TO_EX), .MUX1_SEL(MUX1_SEL), .MUX2_SEL(MUX2_SEL), .UN_SEL(
        UN_SEL), .OP_SEL(OP_SEL), .US_MEM(US_MEM), .TEMP_PC(TEMP_PC), 
        .ALU_OUT({ALU_OUT, EXT_MEM_ADD}), .IMM_OUT(EXT_MEM_DATA), .DEST_OUT(
        DEST_FROM_EXEU) );
  MEMORY_UNIT_NB32_LS5 mem_unit ( .CLK(CLK), .RST(RST), .DEST_IN(
        DEST_FROM_EXEU), .FROM_MEM(EXT_MEM_IN), .FROM_ALU({ALU_OUT, 
        EXT_MEM_ADD}), .ALU_OUT(ALU_TO_WB), .MEM_OUT(TMP_MEM), .DEST_OUT(
        DEST_FROM_MEMU) );
  WRITE_BACK_UNIT_NB32_LS5 wrb_unit ( .MEM_ALU_SEL(MEM_ALU_SEL), .DEST_IN(
        DEST_FROM_MEMU), .FROM_ALU(ALU_TO_WB), .FROM_MEM(TMP_MEM), .DATA_OUT(
        DATA_WB), .DEST_OUT(DEST_FROM_WRBU) );
  FOREWARD_UNIT_NB32_LS5 fw_unit ( .INST_EX({\INST_EX[1] , \INST_EX[0] }), 
        .INST_MEM({\INST_MEM[1] , \INST_MEM[0] }), .INST_T_EX(INST_T_EX), 
        .Rs_EX(RS), .Rt_EX(RT), .Rd_MEM(DEST_FROM_EXEU), .Rd_WB(DEST_FROM_MEMU), .CTL_MUX1(FW_MUX1_SEL), .CTL_MUX2(FW_MUX2_SEL) );
  BUF_X1 U1 ( .A(n6), .Z(FLUSH) );
  INV_X1 U2 ( .A(RST), .ZN(n5) );
  AOI21_X1 U3 ( .B1(MISS_HIT[1]), .B2(MISS_HIT[0]), .A(n5), .ZN(n6) );
endmodule


module DLX ( CLK, RST, D_TYPE, EXT_MEM_IN, IRAM_OUT, RW, US_MEM, IRAM_ADD, 
        EXT_MEM_ADD, EXT_MEM_DATA );
  output [1:0] D_TYPE;
  input [31:0] EXT_MEM_IN;
  input [31:0] IRAM_OUT;
  output [31:0] IRAM_ADD;
  output [4:0] EXT_MEM_ADD;
  output [31:0] EXT_MEM_DATA;
  input CLK, RST;
  output RW, US_MEM;
  wire   STALL, INST_T_EX, JMP, RI, RD1, RD2, WR, PC_SEL, MEM_ALU_SEL, US,
         MUX1_SEL, MUX2_SEL, FLUSH;
  wire   [1:0] INST_EX;
  wire   [1:0] INST_MEM;
  wire   [1:0] BR_TYPE;
  wire   [2:0] UN_SEL;
  wire   [3:0] OP_SEL;
  wire   [10:0] FUNC;
  wire   [5:0] OPCODE;

  DATAPATH_NB32_LS5_OPC6_FN11 dp ( .CLK(CLK), .STALL(STALL), .RST(RST), 
        .INST_EX(INST_EX), .INST_MEM(INST_MEM), .INST_T_EX(INST_T_EX), .JMP(
        JMP), .RI(RI), .RD1(RD1), .RD2(RD2), .WR(WR), .PC_SEL(PC_SEL), 
        .MEM_ALU_SEL(MEM_ALU_SEL), .US(US), .MUX1_SEL(MUX1_SEL), .MUX2_SEL(
        MUX2_SEL), .BR_TYPE(BR_TYPE), .UN_SEL(UN_SEL), .OP_SEL(OP_SEL), 
        .IRAM_OUT(IRAM_OUT), .EXT_MEM_IN(EXT_MEM_IN), .FLUSH(FLUSH), .US_MEM(
        US_MEM), .EXT_MEM_ADD(EXT_MEM_ADD), .EXT_MEM_DATA(EXT_MEM_DATA), 
        .CURR_PC(IRAM_ADD), .FUNC(FUNC), .OP_CODE(OPCODE) );
  DLX_CU cu ( .CLK(CLK), .RST(RST), .OPCODE(OPCODE), .FUNC(FUNC), .FLUSH(FLUSH), .STALL(STALL), .JMP(JMP), .RI(RI), .BR_TYPE(BR_TYPE), .RD1(RD1), .RD2(RD2), 
        .US(US), .MUX1_SEL(MUX1_SEL), .MUX2_SEL(MUX2_SEL), .UN_SEL(UN_SEL), 
        .OP_SEL(OP_SEL), .PC_SEL(PC_SEL), .RW(RW), .D_TYPE(D_TYPE), .WR(WR), 
        .MEM_ALU_SEL(MEM_ALU_SEL), .INST_T_EX(INST_T_EX), .INST_EX(INST_EX), 
        .INST_MEM(INST_MEM) );
endmodule

